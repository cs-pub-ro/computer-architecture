module fpu(
    output wire [31:0] o_w_out,
    input wire [31:0] i_w_op1,
    input wire [31:0] i_w_op2,
    input wire [2:0] i_w_opsel
);

endmodule