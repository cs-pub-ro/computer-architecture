`timescale 1ns / 1ps
module test_mux;
    //Inputs

    //Outputs
    
    //local variables for loop
    integer i,j;

    //Module initialization

    //Simulation tests
    initial begin
        //finish the simulation
        $finish;
    end
endmodule
