module flagram (
    output wire [3:0] o_w_out,
    input wire i_w_clk,
    input wire [3:0] i_w_address,
    input wire [3:0] i_w_data,
    input wire i_w_we,
    input wire i_w_oe,
    input wire i_w_flags_out
);

endmodule
