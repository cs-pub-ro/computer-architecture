module opregister(
    output reg [3:0] o_w_out,
    input wire i_w_clk,
    input wire i_w_reset,
    input wire [3:0] i_w_data,
    input wire i_w_we,
    input wire i_w_oe,
    input wire [1:0] i_w_opsel
);

endmodule