module comb(
    output wire o_w_out,
    input wire i_w_a,
    input wire i_w_b,
    input wire i_w_c
);
    
    //TODO: Implement comb
    assign o_w_out = 1'bz;
endmodule