module led7(
    output wire o_w_ca,
    output wire o_w_cb,
    output wire o_w_cc,
    output wire o_w_cd,
    output wire o_w_ce,
    output wire o_w_cf,
    output wire o_w_cg,
    input wire [1:0] i_w_digit
);

endmodule