module top(input wire [1:0] clock_reset, output wire [15:0] o);
   wire [195:0] od;
   wire [179:0] d;
   wire [217:0] q;
   assign o = od[15:0];
   top_Cu c0(.clock_reset(clock_reset), .i(d[151:125]), .o(q[201:176]));
   top_FR c1(.clock_reset(clock_reset), .i(d[124:109]), .o(q[175:160]));
   top_IR c2(.clock_reset(clock_reset), .i(d[108:93]), .o(q[159:144]));
   top_MA c3(.clock_reset(clock_reset), .i(d[74:57]), .o(q[111:80]));
   top_PC c4(.clock_reset(clock_reset), .i(d[92:75]), .o(q[143:112]));
   top_RAM c5(.clock_reset(clock_reset), .i(d[179:152]), .o(q[217:202]));
   top_T1 c6(.clock_reset(clock_reset), .i(d[38:21]), .o(q[47:16]));
   top_T2 c7(.clock_reset(clock_reset), .i(d[56:39]), .o(q[79:48]));
   top_regs c8(.clock_reset(clock_reset), .i(d[20:0]), .o(q[15:0]));
   assign d = od[195:16];
   assign od = kernel_top_kernel(clock_reset, q);
   function [195:0] kernel_top_kernel(input reg [1:0] arg_0, input reg [217:0] arg_2);
         reg [25:0] or0;
         reg [217:0] or1;
         reg [2:0] or2;
         reg [0:0] or3;
         reg [0:0] or4;
         reg [0:0] or5;
         reg [0:0] or6;
         reg [0:0] or7;
         reg [0:0] or8;
         reg [0:0] or9;
         reg [0:0] or10;
         reg [0:0] or11;
         reg [0:0] or12;
         reg [0:0] or13;
         reg [0:0] or14;
         reg [3:0] or15;
         reg [0:0] or16;
         reg [0:0] or17;
         reg [0:0] or18;
         reg [0:0] or19;
         reg [0:0] or20;
         reg [0:0] or21;
         reg [0:0] or22;
         reg [31:0] or23;
         reg [15:0] or24;
         reg [31:0] or25;
         reg [15:0] or26;
         reg [36:0] or27;
         reg [36:0] or28;
         reg [36:0] or29;
         reg [36:0] or30;
         reg [15:0] or31;
         reg [15:0] or32;
         reg signed [15:0] or33;
         reg [0:0] or34;
         reg signed [15:0] or35;
         reg [0:0] or36;
         reg [0:0] or37;
         reg [0:0] or38;
         reg [15:0] or39;
         reg [3:0] or40;
         reg [16:0] or41;
         reg [16:0] or42;
         reg [16:0] or43;
         reg [17:0] or44;
         reg [17:0] or45;
         reg [17:0] or46;
         reg [1:0] or47;
         reg [17:0] or48;
         reg [0:0] or49;
         // out
         reg [20:0] or50;
         reg [15:0] or51;
         reg [15:0] or52;
         reg [15:0] or53;
         reg [15:0] or54;
         reg [16:0] or55;
         reg [16:0] or56;
         reg [16:0] or57;
         reg [0:0] or58;
         reg [0:0] or59;
         // out
         reg [20:0] or60;
         reg [16:0] or61;
         reg [15:0] or62;
         reg [16:0] or63;
         reg [16:0] or64;
         reg [0:0] or65;
         reg [16:0] or66;
         reg [0:0] or67;
         // out
         reg [20:0] or68;
         reg [15:0] or69;
         reg [0:0] or70;
         reg [0:0] or71;
         // out
         reg [20:0] or72;
         reg [16:0] or73;
         reg [16:0] or74;
         reg signed [16:0] or75;
         reg signed [16:0] or76;
         reg [16:0] or77;
         reg [15:0] or78;
         reg [16:0] or79;
         reg signed [16:0] or80;
         reg [16:0] or81;
         reg [16:0] or82;
         reg [16:0] or83;
         reg signed [16:0] or84;
         reg [0:0] or85;
         // out
         reg [20:0] or86;
         reg signed [16:0] or87;
         reg [16:0] or88;
         reg [15:0] or89;
         reg [16:0] or90;
         reg signed [16:0] or91;
         reg [16:0] or92;
         reg [16:0] or93;
         reg [16:0] or94;
         reg signed [16:0] or95;
         reg [0:0] or96;
         // out
         reg [20:0] or97;
         reg signed [16:0] or98;
         reg [16:0] or99;
         reg [15:0] or100;
         // out
         reg [20:0] or101;
         reg [15:0] or102;
         // out
         reg [20:0] or103;
         reg [15:0] or104;
         reg [0:0] or105;
         reg [0:0] or106;
         // out
         reg [20:0] or107;
         reg [15:0] or108;
         reg signed [15:0] or109;
         reg [0:0] or110;
         // out
         reg [20:0] or111;
         reg [15:0] or112;
         reg [0:0] or113;
         reg [0:0] or114;
         // out
         reg [20:0] or115;
         reg [3:0] or116;
         reg [0:0] or117;
         reg [4:0] or118;
         reg [0:0] or119;
         reg [0:0] or120;
         reg [0:0] or121;
         reg [0:0] or122;
         reg [4:0] or123;
         reg [0:0] or124;
         reg [0:0] or125;
         reg [0:0] or126;
         reg [0:0] or127;
         reg [4:0] or128;
         reg [0:0] or129;
         reg [0:0] or130;
         reg [0:0] or131;
         reg [0:0] or132;
         // out
         reg [20:0] or133;
         reg [15:0] or134;
         reg [15:0] or135;
         reg [15:0] or136;
         reg [7:0] or137;
         reg [15:0] or138;
         reg [7:0] or139;
         reg [15:0] or140;
         reg [15:0] or141;
         reg [15:0] or142;
         reg [31:0] or143;
         reg [15:0] or144;
         reg [15:0] or145;
         reg [15:0] or146;
         reg [15:0] or147;
         reg [15:0] or148;
         reg [15:0] or149;
         reg [15:0] or150;
         reg [15:0] or151;
         reg [15:0] or152;
         reg [17:0] or153;
         reg [17:0] or154;
         reg [17:0] or155;
         // d
         reg [179:0] or156;
         reg [17:0] or157;
         reg [17:0] or158;
         reg [17:0] or159;
         // d
         reg [179:0] or160;
         reg [17:0] or161;
         reg [17:0] or162;
         reg [17:0] or163;
         // d
         reg [179:0] or164;
         reg [31:0] or165;
         reg [15:0] or166;
         reg [9:0] or167;
         reg [27:0] or168;
         reg [27:0] or169;
         reg [27:0] or170;
         reg [27:0] or171;
         // d
         reg [179:0] or172;
         reg [17:0] or173;
         reg [17:0] or174;
         reg [17:0] or175;
         // d
         reg [179:0] or176;
         reg [15:0] or177;
         reg [0:0] or178;
         reg [21:0] or179;
         // d
         reg [179:0] or180;
         reg [15:0] or181;
         reg [0:0] or182;
         reg [0:0] or183;
         reg [14:0] or184;
         reg [15:0] or185;
         reg [0:0] or186;
         reg [0:0] or187;
         reg [13:0] or188;
         reg [15:0] or189;
         reg [0:0] or190;
         reg [0:0] or191;
         reg [12:0] or192;
         reg [15:0] or193;
         reg [0:0] or194;
         reg [0:0] or195;
         reg [11:0] or196;
         reg [15:0] or197;
         reg [0:0] or198;
         reg [0:0] or199;
         reg [4:0] or200;
         reg [4:0] or201;
         reg [4:0] or202;
         reg [4:0] or203;
         reg [4:0] or204;
         // d
         reg [179:0] or205;
         reg [15:0] or206;
         reg [15:0] or207;
         // d
         reg [179:0] or208;
         reg [4:0] or209;
         reg [15:0] or210;
         reg [4:0] or211;
         reg [0:0] or212;
         reg [0:0] or213;
         reg [15:0] or214;
         reg [0:0] or215;
         reg [0:0] or216;
         reg [15:0] or217;
         reg [0:0] or218;
         reg [0:0] or219;
         reg [15:0] or220;
         reg [0:0] or221;
         reg [0:0] or222;
         reg [15:0] or223;
         reg [0:0] or224;
         reg [0:0] or225;
         reg [15:0] or226;
         reg [15:0] or227;
         reg [15:0] or228;
         reg [15:0] or229;
         reg [15:0] or230;
         reg [15:0] or231;
         reg [15:0] or232;
         reg [15:0] or233;
         reg [15:0] or234;
         reg [15:0] or235;
         reg [15:0] or236;
         reg [15:0] or237;
         // d
         reg [179:0] or238;
         reg [17:0] or239;
         reg [17:0] or240;
         reg [17:0] or241;
         // d
         reg [179:0] or242;
         // d
         reg [179:0] or243;
         reg [195:0] or244;
         reg [1:0] or245;
         reg [33:0] or246;
         reg [15:0] or247;
         reg [17:0] or248;
         reg [17:0] or249;
         reg [15:0] or250;
         reg [32:0] or251;
         reg [15:0] or252;
         reg signed [17:0] or253;
         reg [23:0] or254;
         reg [16:0] or255;
         reg [17:0] or256;
         reg [18:0] or257;
         reg [19:0] or258;
         reg [14:0] or259;
         reg [13:0] or260;
         reg [12:0] or261;
         reg [11:0] or262;
         localparam ol0 = 37'b0000000000000000000000000000000000000;
         localparam ol1 = 16'b0000000000000000;
         localparam ol2 = 16'b0000000000000000;
         localparam ol3 = 1'b1;
         localparam ol4 = 1'b0;
         localparam ol5 = 21'bXXXX1XXXXXXXXXXXXXXXX;
         localparam ol6 = 4'b0000;
         localparam ol7 = 4'b0011;
         localparam ol8 = 4'b0100;
         localparam ol9 = 4'b0101;
         localparam ol10 = 4'b0110;
         localparam ol11 = 4'b1000;
         localparam ol12 = 4'b0111;
         localparam ol13 = 4'b1001;
         localparam ol14 = 4'b0001;
         localparam ol15 = 4'b0010;
         localparam ol16 = 16'b0000000000000000;
         localparam ol17 = 4'b0000;
         localparam ol18 = 4'b0001;
         localparam ol19 = 4'b0010;
         localparam ol20 = 1'b0;
         localparam ol21 = 16'b0000000000000000;
         localparam ol22 = 16'b0000000000000000;
         localparam ol23 = 16'b0000000000000000;
         localparam ol24 = 18'b000000000000000000;
         localparam ol25 = 180'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
         localparam ol26 = 18'b000000000000000000;
         localparam ol27 = 18'b000000000000000000;
         localparam ol28 = 28'b0000000000000000000000000000;
         localparam ol29 = 18'b000000000000000000;
         localparam ol30 = 16'b0000000000000000;
         localparam ol31 = 22'b1000000000000000000000;
         localparam ol32 = 22'bXXXXXXXXXXXXXXXXXXXXXX;
         localparam ol33 = 5'b00000;
         localparam ol34 = 1'b1;
         localparam ol35 = 1'b0;
         localparam ol36 = 1'b1;
         localparam ol37 = 1'b0;
         localparam ol38 = 1'b1;
         localparam ol39 = 1'b0;
         localparam ol40 = 1'b1;
         localparam ol41 = 1'b0;
         localparam ol42 = 1'b1;
         localparam ol43 = 1'b0;
         localparam ol44 = 18'b000000000000000000;
         localparam ol45 = 1'b0;
         localparam ol46 = 1'b0;
         localparam ol47 = 1'b0;
         localparam ol48 = 1'b0;
         localparam ol49 = 2'b00;
         localparam ol50 = 3'b000;
         localparam ol51 = 4'b0000;
         begin
            or245 = arg_0;
            or1 = arg_2;
            or0 = or1[201:176];
            or2 = or0[2:0];
            or3 = or0[3:3];
            or4 = or0[4:4];
            or5 = or0[5:5];
            or6 = or0[6:6];
            or7 = or0[7:7];
            or8 = or0[8:8];
            or9 = or0[9:9];
            or10 = or0[10:10];
            or11 = or0[11:11];
            or12 = or0[12:12];
            or13 = or0[13:13];
            or14 = or0[14:14];
            or15 = or0[18:15];
            or16 = or0[19:19];
            or17 = or0[20:20];
            or18 = or0[21:21];
            or19 = or0[22:22];
            or20 = or0[24:24];
            or21 = or0[23:23];
            or22 = or0[25:25];
            or23 = or1[47:16];
            or24 = or23[31:16];
            or25 = or1[79:48];
            or26 = or25[31:16];
            or27 = ol0;
            or27[15:0] = or24;
            or28 = or27;
            or28[31:16] = or26;
            or29 = or28;
            or29[32:32] = or13;
            or30 = or29;
            or30[36:33] = or15;
            or31 = or30[15:0];
            or32 = or30[31:16];
            or33 = $signed(or31);
            or34 = or33 >= ol1;
            or35 = $signed(or32);
            or36 = or35 >= ol2;
            or37 = or30[32:32];
            or38 = or37 ? ol3 : ol4;
            or39 = or31 | or32;
            or40 = or30[36:33];
            or42 = {{1{1'b0}}, or31};
            or43 = {{1{1'b0}}, or32};
            or41 = or42 + or43;
            or45 = {{1{1'b0}}, or41};
            or46 = {{17{1'b0}}, or38};
            or44 = or45 + or46;
            or246 = {{16{1'b0}}, or44};
            or48 = or246[33:16];
            or47 = or48[1:0];
            or49 = |or47;
            or50 = ol5;
            or50[16:16] = or49;
            or51 = or44[15:0];
            or52 = ~or39;
            or53 = or31 & or32;
            or54 = or31 ^ or32;
            or56 = {{1{1'b0}}, or39};
            or247 = or56[15:0];
            or55 = {or247, ol45};
            or248 = {{1{1'b0}}, or55};
            or57 = or248[17:1];
            or58 = or57[0:0];
            or59 = |or58;
            or60 = ol5;
            or60[16:16] = or59;
            or249 = {{1{1'b0}}, or57};
            or61 = or249[17:1];
            or62 = or61[15:0];
            or64 = {{1{1'b0}}, or39};
            or250 = or64[15:0];
            or63 = {or250, ol46};
            or251 = {{16{1'b0}}, or63};
            or66 = or251[32:16];
            or65 = or66[0:0];
            or67 = |or65;
            or68 = ol5;
            or68[16:16] = or67;
            or69 = or63[15:0];
            or70 = or39[0:0];
            or71 = |or70;
            or72 = ol5;
            or72[16:16] = or71;
            or74 = {{1{1'b0}}, or39};
            or252 = or74[15:0];
            or73 = {or252, ol47};
            or75 = $signed(or73);
            or253 = $signed({{1{or75[16]}}, or75});
            or76 = or253[17:1];
            or77 = $unsigned(or76);
            or78 = or77[15:0];
            or79 = {{1{1'b0}}, or31};
            or80 = $signed(or79);
            or82 = {{1{1'b0}}, or32};
            or83 = {{16{1'b0}}, or38};
            or81 = or82 + or83;
            or84 = $signed(or81);
            or85 = or80 > or84;
            or86 = ol5;
            or86[16:16] = or85;
            or87 = or80 - or84;
            or88 = $unsigned(or87);
            or89 = or88[15:0];
            or90 = {{1{1'b0}}, or32};
            or91 = $signed(or90);
            or93 = {{1{1'b0}}, or31};
            or94 = {{16{1'b0}}, or38};
            or92 = or93 + or94;
            or95 = $signed(or92);
            or96 = or91 > or95;
            or97 = ol5;
            or97[16:16] = or96;
            or98 = or91 - or95;
            or99 = $unsigned(or98);
            or100 = or99[15:0];
            case (or40)
               4'b0000 : or101 = or50;
               4'b0011 : or101 = ol5;
               4'b0100 : or101 = ol5;
               4'b0101 : or101 = ol5;
               4'b0110 : or101 = ol5;
               4'b1000 : or101 = or60;
               4'b0111 : or101 = or68;
               4'b1001 : or101 = or72;
               4'b0001 : or101 = or86;
               4'b0010 : or101 = or97;
            endcase
            case (or40)
               4'b0000 : or102 = or51;
               4'b0011 : or102 = or52;
               4'b0100 : or102 = or53;
               4'b0101 : or102 = or39;
               4'b0110 : or102 = or54;
               4'b1000 : or102 = or62;
               4'b0111 : or102 = or69;
               4'b1001 : or102 = or78;
               4'b0001 : or102 = or89;
               4'b0010 : or102 = or100;
            endcase
            or103 = or101;
            or103[15:0] = or102;
            or104 = or103[15:0];
            or105 = |or104;
            or106 = ~or105;
            or107 = or103;
            or107[17:17] = or106;
            or108 = or107[15:0];
            or109 = $signed(or108);
            or110 = or109 < ol16;
            or111 = or107;
            or111[18:18] = or110;
            or112 = or111[15:0];
            or113 = ^or112;
            or114 = ~or113;
            or115 = or111;
            or115[20:20] = or114;
            or116 = or30[36:33];
            or117 = or34 == or36;
            or118 = or115[20:16];
            or119 = or118[2:2];
            or120 = or34 != or119;
            or121 = or117 & or120;
            or122 = or34 != or36;
            or123 = or115[20:16];
            or124 = or123[2:2];
            or125 = or34 != or124;
            or126 = or122 & or125;
            or127 = or36 != or34;
            or128 = or115[20:16];
            or129 = or128[2:2];
            or130 = or36 != or129;
            or131 = or127 & or130;
            case (or116)
               4'b0000 : or132 = or121;
               4'b0001 : or132 = or126;
               4'b0010 : or132 = or131;
               default : or132 = ol20;
            endcase
            or133 = or115;
            or133[19:19] = or132;
            or134 = or1[175:160];
            or135 = or20 ? or134 : ol21;
            or136 = or1[159:144];
            or254 = {{8{1'b0}}, or136};
            or138 = or254[23:8];
            or137 = or138[7:0];
            or139 = or137[7:0];
            or140 = {{8{1'b0}}, or139};
            or141 = or19 ? or140 : ol22;
            or142 = or135 | or141;
            or143 = or1[143:112];
            or144 = or143[15:0];
            or145 = or142 | or144;
            or146 = or1[15:0];
            or147 = or145 | or146;
            or148 = or1[217:202];
            or149 = or147 | or148;
            or150 = or133[15:0];
            or151 = or14 ? or150 : ol23;
            or152 = or149 | or151;
            or153 = ol24;
            or153[16:16] = or5;
            or154 = or153;
            or154[17:17] = or6;
            or155 = or154;
            or155[15:0] = or152;
            or156 = ol25;
            or156[38:21] = or155;
            or157 = ol26;
            or157[16:16] = or7;
            or158 = or157;
            or158[17:17] = or8;
            or159 = or158;
            or159[15:0] = or152;
            or160 = or156;
            or160[56:39] = or159;
            or161 = ol27;
            or161[16:16] = or9;
            or162 = or161;
            or162[17:17] = or10;
            or163 = or162;
            or163[15:0] = or152;
            or164 = or160;
            or164[74:57] = or163;
            or165 = or1[111:80];
            or166 = or165[31:16];
            or167 = or166[9:0];
            or168 = ol28;
            or168[0:0] = or11;
            or169 = or168;
            or169[1:1] = or12;
            or170 = or169;
            or170[17:2] = or152;
            or171 = or170;
            or171[27:18] = or167;
            or172 = or164;
            or172[179:152] = or171;
            or173 = ol29;
            or173[15:0] = or152;
            or174 = or173;
            or174[16:16] = or17;
            or175 = or174;
            or175[17:17] = or16;
            or176 = or172;
            or176[92:75] = or175;
            or177 = or1[159:144];
            or178 = or177 == ol30;
            or179 = or178 ? ol31 : ol32;
            or180 = or176;
            or180[146:125] = or179;
            or181 = or1[175:160];
            or182 = or181[0:0];
            or183 = |or182;
            or255 = {{1{1'b0}}, or181};
            or185 = or255[16:1];
            or184 = or185[14:0];
            or186 = or184[0:0];
            or187 = |or186;
            or256 = {{2{1'b0}}, or181};
            or189 = or256[17:2];
            or188 = or189[13:0];
            or190 = or188[0:0];
            or191 = |or190;
            or257 = {{3{1'b0}}, or181};
            or193 = or257[18:3];
            or192 = or193[12:0];
            or194 = or192[0:0];
            or195 = |or194;
            or258 = {{4{1'b0}}, or181};
            or197 = or258[19:4];
            or196 = or197[11:0];
            or198 = or196[0:0];
            or199 = |or198;
            or200 = ol33;
            or200[0:0] = or183;
            or201 = or200;
            or201[1:1] = or187;
            or202 = or201;
            or202[2:2] = or191;
            or203 = or202;
            or203[3:3] = or195;
            or204 = or203;
            or204[4:4] = or199;
            or205 = or180;
            or205[151:147] = or204;
            or206 = or1[159:144];
            or207 = or18 ? or152 : or206;
            or208 = or205;
            or208[108:93] = or207;
            or209 = or152[4:0];
            or210 = {{11{1'b0}}, or209};
            or211 = or133[20:16];
            or212 = or211[0:0];
            or213 = or212 ? ol34 : ol35;
            or214 = {{15{1'b0}}, or213};
            or215 = or211[1:1];
            or216 = or215 ? ol36 : ol37;
            or217 = {{15{1'b0}}, or216};
            or218 = or211[2:2];
            or219 = or218 ? ol38 : ol39;
            or220 = {{15{1'b0}}, or219};
            or221 = or211[3:3];
            or222 = or221 ? ol40 : ol41;
            or223 = {{15{1'b0}}, or222};
            or224 = or211[4:4];
            or225 = or224 ? ol42 : ol43;
            or226 = {{15{1'b0}}, or225};
            or259 = or217[14:0];
            or227 = {or259, ol48};
            or228 = or214 | or227;
            or260 = or220[13:0];
            or229 = {or260, ol49};
            or230 = or228 | or229;
            or261 = or223[12:0];
            or231 = {or261, ol50};
            or232 = or230 | or231;
            or262 = or226[11:0];
            or233 = {or262, ol51};
            or234 = or232 | or233;
            or235 = or22 ? or210 : or234;
            or236 = or1[175:160];
            or237 = or21 ? or235 : or236;
            or238 = or208;
            or238[124:109] = or237;
            or239 = ol44;
            or239[16:16] = or3;
            or240 = or239;
            or240[17:17] = or4;
            or241 = or240;
            or241[15:0] = or152;
            or242 = or238;
            or242[17:0] = or241;
            or243 = or242;
            or243[20:18] = or2;
            or244 = {or243, or152};
            kernel_top_kernel = or244;
         end
   endfunction
endmodule
module top_Cu(input wire [1:0] clock_reset, input wire [26:0] i, output wire [25:0] o);
   wire [28:0] od;
   wire [2:0] d;
   wire [2:0] q;
   assign o = od[25:0];
   top_Cu_state c0(.clock_reset(clock_reset), .i(d[2:0]), .o(q[2:0]));
   assign d = od[28:26];
   assign od = kernel_cu_kernel(clock_reset, i, q);
   function [28:0] kernel_cu_kernel(input reg [1:0] arg_0, input reg [26:0] arg_1, input reg [2:0] arg_2);
         reg [2:0] or0;
         // cs
         reg [25:0] or1;
         reg [2:0] or2;
         reg [2:0] or3;
         reg [28:0] or4;
         reg [1:0] or5;
         reg [26:0] or6;
         localparam ol0 = 3'b000;
         localparam ol1 = 26'b00000000000000000000000000;
         localparam ol2 = 3'b001;
         localparam ol3 = 3'b010;
         localparam ol4 = 3'b011;
         localparam ol5 = 3'b100;
         localparam ol6 = 3'b101;
         localparam ol7 = 26'b00000100000000000001000000;
         localparam ol8 = 3'b110;
         localparam ol9 = 26'b00000010000110000000100000;
         localparam ol10 = 3'b111;
         localparam ol11 = 3'b001;
         localparam ol12 = 3'b010;
         localparam ol13 = 3'b011;
         localparam ol14 = 3'b100;
         localparam ol15 = 3'b101;
         localparam ol16 = 3'b110;
         localparam ol17 = 3'b001;
         localparam ol18 = 3'b111;
         localparam ol19 = 3'b000;
         begin
            or5 = arg_0;
            or6 = arg_1;
            or0 = arg_2;
            case (or0)
               3'b000 : or1 = ol1;
               3'b001 : or1 = ol1;
               3'b010 : or1 = ol1;
               3'b011 : or1 = ol1;
               3'b100 : or1 = ol1;
               3'b101 : or1 = ol7;
               3'b110 : or1 = ol9;
               3'b111 : or1 = ol1;
            endcase
            case (or0)
               3'b000 : or2 = ol11;
               3'b001 : or2 = ol12;
               3'b010 : or2 = ol13;
               3'b011 : or2 = ol14;
               3'b100 : or2 = ol15;
               3'b101 : or2 = ol16;
               3'b110 : or2 = ol17;
               3'b111 : or2 = ol18;
            endcase
            or3 = ol19;
            or3[2:0] = or2;
            or4 = {or3, or1};
            kernel_cu_kernel = or4;
         end
   endfunction
endmodule
module top_Cu_state(input wire [1:0] clock_reset, input wire [2:0] i, output reg [2:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 3'b000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 3'b000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_FR(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_IR(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_MA(input wire [1:0] clock_reset, input wire [17:0] i, output wire [31:0] o);
   wire [47:0] od;
   wire [15:0] d;
   wire [15:0] q;
   assign o = od[31:0];
   top_MA_memory c0(.clock_reset(clock_reset), .i(d[15:0]), .o(q[15:0]));
   assign d = od[47:32];
   assign od = kernel_reg_ker(clock_reset, i, q);
   function [47:0] kernel_reg_ker(input reg [1:0] arg_0, input reg [17:0] arg_1, input reg [15:0] arg_2);
         reg [0:0] or0;
         reg [17:0] or1;
         reg [0:0] or2;
         reg [0:0] or3;
         reg [0:0] or4;
         reg [15:0] or5;
         reg [15:0] or6;
         reg [0:0] or7;
         reg [15:0] or8;
         reg [31:0] or9;
         reg [0:0] or10;
         reg [15:0] or11;
         reg [15:0] or12;
         reg [15:0] or13;
         reg [47:0] or14;
         reg [1:0] or15;
         localparam ol0 = 16'b0000000000000000;
         localparam ol1 = 16'b0000000000000000;
         localparam ol2 = 16'b0000000000000000;
         begin
            or15 = arg_0;
            or1 = arg_1;
            or5 = arg_2;
            or0 = or1[16:16];
            or2 = or1[17:17];
            or3 = ~or2;
            or4 = or0 & or3;
            or6 = or4 ? or5 : ol0;
            or7 = or1[16:16];
            or8 = or7 ? or5 : ol1;
            or9 = {or8, or6};
            or10 = or1[17:17];
            or11 = or1[15:0];
            or12 = or10 ? or11 : or5;
            or13 = ol2;
            or13[15:0] = or12;
            or14 = {or13, or9};
            kernel_reg_ker = or14;
         end
   endfunction
endmodule
module top_MA_memory(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_PC(input wire [1:0] clock_reset, input wire [17:0] i, output wire [31:0] o);
   wire [47:0] od;
   wire [15:0] d;
   wire [15:0] q;
   assign o = od[31:0];
   top_PC_memory c0(.clock_reset(clock_reset), .i(d[15:0]), .o(q[15:0]));
   assign d = od[47:32];
   assign od = kernel_reg_ker(clock_reset, i, q);
   function [47:0] kernel_reg_ker(input reg [1:0] arg_0, input reg [17:0] arg_1, input reg [15:0] arg_2);
         reg [0:0] or0;
         reg [17:0] or1;
         reg [0:0] or2;
         reg [0:0] or3;
         reg [0:0] or4;
         reg [15:0] or5;
         reg [15:0] or6;
         reg [0:0] or7;
         reg [15:0] or8;
         reg [31:0] or9;
         reg [0:0] or10;
         reg [15:0] or11;
         reg [15:0] or12;
         reg [15:0] or13;
         reg [47:0] or14;
         reg [1:0] or15;
         localparam ol0 = 16'b0000000000000000;
         localparam ol1 = 16'b0000000000000000;
         localparam ol2 = 16'b0000000000000000;
         begin
            or15 = arg_0;
            or1 = arg_1;
            or5 = arg_2;
            or0 = or1[16:16];
            or2 = or1[17:17];
            or3 = ~or2;
            or4 = or0 & or3;
            or6 = or4 ? or5 : ol0;
            or7 = or1[16:16];
            or8 = or7 ? or5 : ol1;
            or9 = {or8, or6};
            or10 = or1[17:17];
            or11 = or1[15:0];
            or12 = or10 ? or11 : or5;
            or13 = ol2;
            or13[15:0] = or12;
            or14 = {or13, or9};
            kernel_reg_ker = or14;
         end
   endfunction
endmodule
module top_PC_memory(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_RAM(input wire [1:0] clock_reset, input wire [27:0] i, output wire [15:0] o);
   wire [52:0] od;
   wire [36:0] d;
   wire [15:0] q;
   assign o = od[15:0];
   top_RAM_memory c0(.clock_reset(clock_reset), .i(d[36:0]), .o(q[15:0]));
   assign d = od[52:16];
   assign od = kernel_ram_kernel(clock_reset, i, q);
   function [52:0] kernel_ram_kernel(input reg [1:0] arg_0, input reg [27:0] arg_1, input reg [15:0] arg_2);
         reg [9:0] or0;
         reg [27:0] or1;
         // d
         reg [36:0] or2;
         reg [9:0] or3;
         reg [15:0] or4;
         reg [0:0] or5;
         reg [26:0] or6;
         reg [26:0] or7;
         reg [26:0] or8;
         // d
         reg [36:0] or9;
         reg [0:0] or10;
         reg [0:0] or11;
         reg [0:0] or12;
         reg [0:0] or13;
         reg [15:0] or14;
         reg [15:0] or15;
         reg [52:0] or16;
         reg [1:0] or17;
         localparam ol0 = 37'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
         localparam ol1 = 27'b000000000000000000000000000;
         localparam ol2 = 16'b0000000000000000;
         begin
            or17 = arg_0;
            or1 = arg_1;
            or14 = arg_2;
            or0 = or1[27:18];
            or2 = ol0;
            or2[9:0] = or0;
            or3 = or1[27:18];
            or4 = or1[17:2];
            or5 = or1[1:1];
            or6 = ol1;
            or6[9:0] = or3;
            or7 = or6;
            or7[25:10] = or4;
            or8 = or7;
            or8[26:26] = or5;
            or9 = or2;
            or9[36:10] = or8;
            or10 = or1[0:0];
            or11 = or1[1:1];
            or12 = ~or11;
            or13 = or10 & or12;
            or15 = or13 ? or14 : ol2;
            or16 = {or9, or15};
            kernel_ram_kernel = or16;
         end
   endfunction
endmodule
module top_RAM_memory(input wire [1:0] clock_reset, input wire [36:0] i, output reg [15:0] o);
   wire [9:0] read_addr;
   wire [9:0] write_addr;
   wire [15:0] write_value;
   wire [0:0] write_enable;
   wire [0:0] clock;
   reg [15:0] mem[1023:0];
   initial begin
      mem[0] = 16'b0000000000110001;
      mem[1] = 16'b0100001010010010;
      mem[2] = 16'b0110000100101110;
      mem[3] = 16'b0000000000101011;
      mem[4] = 16'b0000000000101010;
      mem[5] = 16'b0000001100001000;
      mem[6] = 16'b1110000000001000;
      mem[7] = 16'b0110001000001000;
      mem[8] = 16'b0000000000101011;
      mem[9] = 16'b1110001000001000;
      mem[10] = 16'b0000000000001100;
      mem[11] = 16'b0010000100001000;
      mem[12] = 16'b0000000000010111;
      mem[13] = 16'b0110000100001000;
      mem[14] = 16'b0000000000101010;
      mem[15] = 16'b1110000100001000;
      mem[16] = 16'b0000000000000001;
      mem[17] = 16'b1100000000001000;
      mem[18] = 16'b0100000000001000;
      mem[19] = 16'b0100000000001000;
      mem[20] = 16'b1100001000001000;
      mem[21] = 16'b1010001000001000;
      mem[22] = 16'b1100000100001000;
      mem[23] = 16'b0000000000000010;
      mem[24] = 16'b0000000000000000;
      mem[25] = 16'b0000000000000000;
      mem[26] = 16'b0000000000000000;
      mem[27] = 16'b0000000000000000;
      mem[28] = 16'b0000000000000000;
      mem[29] = 16'b0000000000000000;
      mem[30] = 16'b0000000000000000;
      mem[31] = 16'b0000000000000000;
      mem[32] = 16'b0000000000000000;
      mem[33] = 16'b0000000000000000;
      mem[34] = 16'b0000000000000000;
      mem[35] = 16'b0000000000000000;
      mem[36] = 16'b0000000000000000;
      mem[37] = 16'b0000000000000000;
      mem[38] = 16'b0000000000000000;
      mem[39] = 16'b0000000000000000;
      mem[40] = 16'b0000000000000000;
      mem[41] = 16'b0000000000000000;
      mem[42] = 16'b0000000000000000;
      mem[43] = 16'b0000000000000000;
      mem[44] = 16'b0000000000000000;
      mem[45] = 16'b0000000000000000;
      mem[46] = 16'b0000000000000000;
      mem[47] = 16'b0000000000000000;
      mem[48] = 16'b0000000000000000;
      mem[49] = 16'b0000000000000000;
      mem[50] = 16'b0000000000000000;
      mem[51] = 16'b0000000000000000;
      mem[52] = 16'b0000000000000000;
      mem[53] = 16'b0000000000000000;
      mem[54] = 16'b0000000000000000;
      mem[55] = 16'b0000000000000000;
      mem[56] = 16'b0000000000000000;
      mem[57] = 16'b0000000000000000;
      mem[58] = 16'b0000000000000000;
      mem[59] = 16'b0000000000000000;
      mem[60] = 16'b0000000000000000;
      mem[61] = 16'b0000000000000000;
      mem[62] = 16'b0000000000000000;
      mem[63] = 16'b0000000000000000;
      mem[64] = 16'b0000000000000000;
      mem[65] = 16'b0000000000000000;
      mem[66] = 16'b0000000000000000;
      mem[67] = 16'b0000000000000000;
      mem[68] = 16'b0000000000000000;
      mem[69] = 16'b0000000000000000;
      mem[70] = 16'b0000000000000000;
      mem[71] = 16'b0000000000000000;
      mem[72] = 16'b0000000000000000;
      mem[73] = 16'b0000000000000000;
      mem[74] = 16'b0000000000000000;
      mem[75] = 16'b0000000000000000;
      mem[76] = 16'b0000000000000000;
      mem[77] = 16'b0000000000000000;
      mem[78] = 16'b0000000000000000;
      mem[79] = 16'b0000000000000000;
      mem[80] = 16'b0000000000000000;
      mem[81] = 16'b0000000000000000;
      mem[82] = 16'b0000000000000000;
      mem[83] = 16'b0000000000000000;
      mem[84] = 16'b0000000000000000;
      mem[85] = 16'b0000000000000000;
      mem[86] = 16'b0000000000000000;
      mem[87] = 16'b0000000000000000;
      mem[88] = 16'b0000000000000000;
      mem[89] = 16'b0000000000000000;
      mem[90] = 16'b0000000000000000;
      mem[91] = 16'b0000000000000000;
      mem[92] = 16'b0000000000000000;
      mem[93] = 16'b0000000000000000;
      mem[94] = 16'b0000000000000000;
      mem[95] = 16'b0000000000000000;
      mem[96] = 16'b0000000000000000;
      mem[97] = 16'b0000000000000000;
      mem[98] = 16'b0000000000000000;
      mem[99] = 16'b0000000000000000;
      mem[100] = 16'b0000000000000000;
      mem[101] = 16'b0000000000000000;
      mem[102] = 16'b0000000000000000;
      mem[103] = 16'b0000000000000000;
      mem[104] = 16'b0000000000000000;
      mem[105] = 16'b0000000000000000;
      mem[106] = 16'b0000000000000000;
      mem[107] = 16'b0000000000000000;
      mem[108] = 16'b0000000000000000;
      mem[109] = 16'b0000000000000000;
      mem[110] = 16'b0000000000000000;
      mem[111] = 16'b0000000000000000;
      mem[112] = 16'b0000000000000000;
      mem[113] = 16'b0000000000000000;
      mem[114] = 16'b0000000000000000;
      mem[115] = 16'b0000000000000000;
      mem[116] = 16'b0000000000000000;
      mem[117] = 16'b0000000000000000;
      mem[118] = 16'b0000000000000000;
      mem[119] = 16'b0000000000000000;
      mem[120] = 16'b0000000000000000;
      mem[121] = 16'b0000000000000000;
      mem[122] = 16'b0000000000000000;
      mem[123] = 16'b0000000000000000;
      mem[124] = 16'b0000000000000000;
      mem[125] = 16'b0000000000000000;
      mem[126] = 16'b0000000000000000;
      mem[127] = 16'b0000000000000000;
      mem[128] = 16'b0000000000000000;
      mem[129] = 16'b0000000000000000;
      mem[130] = 16'b0000000000000000;
      mem[131] = 16'b0000000000000000;
      mem[132] = 16'b0000000000000000;
      mem[133] = 16'b0000000000000000;
      mem[134] = 16'b0000000000000000;
      mem[135] = 16'b0000000000000000;
      mem[136] = 16'b0000000000000000;
      mem[137] = 16'b0000000000000000;
      mem[138] = 16'b0000000000000000;
      mem[139] = 16'b0000000000000000;
      mem[140] = 16'b0000000000000000;
      mem[141] = 16'b0000000000000000;
      mem[142] = 16'b0000000000000000;
      mem[143] = 16'b0000000000000000;
      mem[144] = 16'b0000000000000000;
      mem[145] = 16'b0000000000000000;
      mem[146] = 16'b0000000000000000;
      mem[147] = 16'b0000000000000000;
      mem[148] = 16'b0000000000000000;
      mem[149] = 16'b0000000000000000;
      mem[150] = 16'b0000000000000000;
      mem[151] = 16'b0000000000000000;
      mem[152] = 16'b0000000000000000;
      mem[153] = 16'b0000000000000000;
      mem[154] = 16'b0000000000000000;
      mem[155] = 16'b0000000000000000;
      mem[156] = 16'b0000000000000000;
      mem[157] = 16'b0000000000000000;
      mem[158] = 16'b0000000000000000;
      mem[159] = 16'b0000000000000000;
      mem[160] = 16'b0000000000000000;
      mem[161] = 16'b0000000000000000;
      mem[162] = 16'b0000000000000000;
      mem[163] = 16'b0000000000000000;
      mem[164] = 16'b0000000000000000;
      mem[165] = 16'b0000000000000000;
      mem[166] = 16'b0000000000000000;
      mem[167] = 16'b0000000000000000;
      mem[168] = 16'b0000000000000000;
      mem[169] = 16'b0000000000000000;
      mem[170] = 16'b0000000000000000;
      mem[171] = 16'b0000000000000000;
      mem[172] = 16'b0000000000000000;
      mem[173] = 16'b0000000000000000;
      mem[174] = 16'b0000000000000000;
      mem[175] = 16'b0000000000000000;
      mem[176] = 16'b0000000000000000;
      mem[177] = 16'b0000000000000000;
      mem[178] = 16'b0000000000000000;
      mem[179] = 16'b0000000000000000;
      mem[180] = 16'b0000000000000000;
      mem[181] = 16'b0000000000000000;
      mem[182] = 16'b0000000000000000;
      mem[183] = 16'b0000000000000000;
      mem[184] = 16'b0000000000000000;
      mem[185] = 16'b0000000000000000;
      mem[186] = 16'b0000000000000000;
      mem[187] = 16'b0000000000000000;
      mem[188] = 16'b0000000000000000;
      mem[189] = 16'b0000000000000000;
      mem[190] = 16'b0000000000000000;
      mem[191] = 16'b0000000000000000;
      mem[192] = 16'b0000000000000000;
      mem[193] = 16'b0000000000000000;
      mem[194] = 16'b0000000000000000;
      mem[195] = 16'b0000000000000000;
      mem[196] = 16'b0000000000000000;
      mem[197] = 16'b0000000000000000;
      mem[198] = 16'b0000000000000000;
      mem[199] = 16'b0000000000000000;
      mem[200] = 16'b0000000000000000;
      mem[201] = 16'b0000000000000000;
      mem[202] = 16'b0000000000000000;
      mem[203] = 16'b0000000000000000;
      mem[204] = 16'b0000000000000000;
      mem[205] = 16'b0000000000000000;
      mem[206] = 16'b0000000000000000;
      mem[207] = 16'b0000000000000000;
      mem[208] = 16'b0000000000000000;
      mem[209] = 16'b0000000000000000;
      mem[210] = 16'b0000000000000000;
      mem[211] = 16'b0000000000000000;
      mem[212] = 16'b0000000000000000;
      mem[213] = 16'b0000000000000000;
      mem[214] = 16'b0000000000000000;
      mem[215] = 16'b0000000000000000;
      mem[216] = 16'b0000000000000000;
      mem[217] = 16'b0000000000000000;
      mem[218] = 16'b0000000000000000;
      mem[219] = 16'b0000000000000000;
      mem[220] = 16'b0000000000000000;
      mem[221] = 16'b0000000000000000;
      mem[222] = 16'b0000000000000000;
      mem[223] = 16'b0000000000000000;
      mem[224] = 16'b0000000000000000;
      mem[225] = 16'b0000000000000000;
      mem[226] = 16'b0000000000000000;
      mem[227] = 16'b0000000000000000;
      mem[228] = 16'b0000000000000000;
      mem[229] = 16'b0000000000000000;
      mem[230] = 16'b0000000000000000;
      mem[231] = 16'b0000000000000000;
      mem[232] = 16'b0000000000000000;
      mem[233] = 16'b0000000000000000;
      mem[234] = 16'b0000000000000000;
      mem[235] = 16'b0000000000000000;
      mem[236] = 16'b0000000000000000;
      mem[237] = 16'b0000000000000000;
      mem[238] = 16'b0000000000000000;
      mem[239] = 16'b0000000000000000;
      mem[240] = 16'b0000000000000000;
      mem[241] = 16'b0000000000000000;
      mem[242] = 16'b0000000000000000;
      mem[243] = 16'b0000000000000000;
      mem[244] = 16'b0000000000000000;
      mem[245] = 16'b0000000000000000;
      mem[246] = 16'b0000000000000000;
      mem[247] = 16'b0000000000000000;
      mem[248] = 16'b0000000000000000;
      mem[249] = 16'b0000000000000000;
      mem[250] = 16'b0000000000000000;
      mem[251] = 16'b0000000000000000;
      mem[252] = 16'b0000000000000000;
      mem[253] = 16'b0000000000000000;
      mem[254] = 16'b0000000000000000;
      mem[255] = 16'b0000000000000000;
      mem[256] = 16'b0000000000000000;
      mem[257] = 16'b0000000000000000;
      mem[258] = 16'b0000000000000000;
      mem[259] = 16'b0000000000000000;
      mem[260] = 16'b0000000000000000;
      mem[261] = 16'b0000000000000000;
      mem[262] = 16'b0000000000000000;
      mem[263] = 16'b0000000000000000;
      mem[264] = 16'b0000000000000000;
      mem[265] = 16'b0000000000000000;
      mem[266] = 16'b0000000000000000;
      mem[267] = 16'b0000000000000000;
      mem[268] = 16'b0000000000000000;
      mem[269] = 16'b0000000000000000;
      mem[270] = 16'b0000000000000000;
      mem[271] = 16'b0000000000000000;
      mem[272] = 16'b0000000000000000;
      mem[273] = 16'b0000000000000000;
      mem[274] = 16'b0000000000000000;
      mem[275] = 16'b0000000000000000;
      mem[276] = 16'b0000000000000000;
      mem[277] = 16'b0000000000000000;
      mem[278] = 16'b0000000000000000;
      mem[279] = 16'b0000000000000000;
      mem[280] = 16'b0000000000000000;
      mem[281] = 16'b0000000000000000;
      mem[282] = 16'b0000000000000000;
      mem[283] = 16'b0000000000000000;
      mem[284] = 16'b0000000000000000;
      mem[285] = 16'b0000000000000000;
      mem[286] = 16'b0000000000000000;
      mem[287] = 16'b0000000000000000;
      mem[288] = 16'b0000000000000000;
      mem[289] = 16'b0000000000000000;
      mem[290] = 16'b0000000000000000;
      mem[291] = 16'b0000000000000000;
      mem[292] = 16'b0000000000000000;
      mem[293] = 16'b0000000000000000;
      mem[294] = 16'b0000000000000000;
      mem[295] = 16'b0000000000000000;
      mem[296] = 16'b0000000000000000;
      mem[297] = 16'b0000000000000000;
      mem[298] = 16'b0000000000000000;
      mem[299] = 16'b0000000000000000;
      mem[300] = 16'b0000000000000000;
      mem[301] = 16'b0000000000000000;
      mem[302] = 16'b0000000000000000;
      mem[303] = 16'b0000000000000000;
      mem[304] = 16'b0000000000000000;
      mem[305] = 16'b0000000000000000;
      mem[306] = 16'b0000000000000000;
      mem[307] = 16'b0000000000000000;
      mem[308] = 16'b0000000000000000;
      mem[309] = 16'b0000000000000000;
      mem[310] = 16'b0000000000000000;
      mem[311] = 16'b0000000000000000;
      mem[312] = 16'b0000000000000000;
      mem[313] = 16'b0000000000000000;
      mem[314] = 16'b0000000000000000;
      mem[315] = 16'b0000000000000000;
      mem[316] = 16'b0000000000000000;
      mem[317] = 16'b0000000000000000;
      mem[318] = 16'b0000000000000000;
      mem[319] = 16'b0000000000000000;
      mem[320] = 16'b0000000000000000;
      mem[321] = 16'b0000000000000000;
      mem[322] = 16'b0000000000000000;
      mem[323] = 16'b0000000000000000;
      mem[324] = 16'b0000000000000000;
      mem[325] = 16'b0000000000000000;
      mem[326] = 16'b0000000000000000;
      mem[327] = 16'b0000000000000000;
      mem[328] = 16'b0000000000000000;
      mem[329] = 16'b0000000000000000;
      mem[330] = 16'b0000000000000000;
      mem[331] = 16'b0000000000000000;
      mem[332] = 16'b0000000000000000;
      mem[333] = 16'b0000000000000000;
      mem[334] = 16'b0000000000000000;
      mem[335] = 16'b0000000000000000;
      mem[336] = 16'b0000000000000000;
      mem[337] = 16'b0000000000000000;
      mem[338] = 16'b0000000000000000;
      mem[339] = 16'b0000000000000000;
      mem[340] = 16'b0000000000000000;
      mem[341] = 16'b0000000000000000;
      mem[342] = 16'b0000000000000000;
      mem[343] = 16'b0000000000000000;
      mem[344] = 16'b0000000000000000;
      mem[345] = 16'b0000000000000000;
      mem[346] = 16'b0000000000000000;
      mem[347] = 16'b0000000000000000;
      mem[348] = 16'b0000000000000000;
      mem[349] = 16'b0000000000000000;
      mem[350] = 16'b0000000000000000;
      mem[351] = 16'b0000000000000000;
      mem[352] = 16'b0000000000000000;
      mem[353] = 16'b0000000000000000;
      mem[354] = 16'b0000000000000000;
      mem[355] = 16'b0000000000000000;
      mem[356] = 16'b0000000000000000;
      mem[357] = 16'b0000000000000000;
      mem[358] = 16'b0000000000000000;
      mem[359] = 16'b0000000000000000;
      mem[360] = 16'b0000000000000000;
      mem[361] = 16'b0000000000000000;
      mem[362] = 16'b0000000000000000;
      mem[363] = 16'b0000000000000000;
      mem[364] = 16'b0000000000000000;
      mem[365] = 16'b0000000000000000;
      mem[366] = 16'b0000000000000000;
      mem[367] = 16'b0000000000000000;
      mem[368] = 16'b0000000000000000;
      mem[369] = 16'b0000000000000000;
      mem[370] = 16'b0000000000000000;
      mem[371] = 16'b0000000000000000;
      mem[372] = 16'b0000000000000000;
      mem[373] = 16'b0000000000000000;
      mem[374] = 16'b0000000000000000;
      mem[375] = 16'b0000000000000000;
      mem[376] = 16'b0000000000000000;
      mem[377] = 16'b0000000000000000;
      mem[378] = 16'b0000000000000000;
      mem[379] = 16'b0000000000000000;
      mem[380] = 16'b0000000000000000;
      mem[381] = 16'b0000000000000000;
      mem[382] = 16'b0000000000000000;
      mem[383] = 16'b0000000000000000;
      mem[384] = 16'b0000000000000000;
      mem[385] = 16'b0000000000000000;
      mem[386] = 16'b0000000000000000;
      mem[387] = 16'b0000000000000000;
      mem[388] = 16'b0000000000000000;
      mem[389] = 16'b0000000000000000;
      mem[390] = 16'b0000000000000000;
      mem[391] = 16'b0000000000000000;
      mem[392] = 16'b0000000000000000;
      mem[393] = 16'b0000000000000000;
      mem[394] = 16'b0000000000000000;
      mem[395] = 16'b0000000000000000;
      mem[396] = 16'b0000000000000000;
      mem[397] = 16'b0000000000000000;
      mem[398] = 16'b0000000000000000;
      mem[399] = 16'b0000000000000000;
      mem[400] = 16'b0000000000000000;
      mem[401] = 16'b0000000000000000;
      mem[402] = 16'b0000000000000000;
      mem[403] = 16'b0000000000000000;
      mem[404] = 16'b0000000000000000;
      mem[405] = 16'b0000000000000000;
      mem[406] = 16'b0000000000000000;
      mem[407] = 16'b0000000000000000;
      mem[408] = 16'b0000000000000000;
      mem[409] = 16'b0000000000000000;
      mem[410] = 16'b0000000000000000;
      mem[411] = 16'b0000000000000000;
      mem[412] = 16'b0000000000000000;
      mem[413] = 16'b0000000000000000;
      mem[414] = 16'b0000000000000000;
      mem[415] = 16'b0000000000000000;
      mem[416] = 16'b0000000000000000;
      mem[417] = 16'b0000000000000000;
      mem[418] = 16'b0000000000000000;
      mem[419] = 16'b0000000000000000;
      mem[420] = 16'b0000000000000000;
      mem[421] = 16'b0000000000000000;
      mem[422] = 16'b0000000000000000;
      mem[423] = 16'b0000000000000000;
      mem[424] = 16'b0000000000000000;
      mem[425] = 16'b0000000000000000;
      mem[426] = 16'b0000000000000000;
      mem[427] = 16'b0000000000000000;
      mem[428] = 16'b0000000000000000;
      mem[429] = 16'b0000000000000000;
      mem[430] = 16'b0000000000000000;
      mem[431] = 16'b0000000000000000;
      mem[432] = 16'b0000000000000000;
      mem[433] = 16'b0000000000000000;
      mem[434] = 16'b0000000000000000;
      mem[435] = 16'b0000000000000000;
      mem[436] = 16'b0000000000000000;
      mem[437] = 16'b0000000000000000;
      mem[438] = 16'b0000000000000000;
      mem[439] = 16'b0000000000000000;
      mem[440] = 16'b0000000000000000;
      mem[441] = 16'b0000000000000000;
      mem[442] = 16'b0000000000000000;
      mem[443] = 16'b0000000000000000;
      mem[444] = 16'b0000000000000000;
      mem[445] = 16'b0000000000000000;
      mem[446] = 16'b0000000000000000;
      mem[447] = 16'b0000000000000000;
      mem[448] = 16'b0000000000000000;
      mem[449] = 16'b0000000000000000;
      mem[450] = 16'b0000000000000000;
      mem[451] = 16'b0000000000000000;
      mem[452] = 16'b0000000000000000;
      mem[453] = 16'b0000000000000000;
      mem[454] = 16'b0000000000000000;
      mem[455] = 16'b0000000000000000;
      mem[456] = 16'b0000000000000000;
      mem[457] = 16'b0000000000000000;
      mem[458] = 16'b0000000000000000;
      mem[459] = 16'b0000000000000000;
      mem[460] = 16'b0000000000000000;
      mem[461] = 16'b0000000000000000;
      mem[462] = 16'b0000000000000000;
      mem[463] = 16'b0000000000000000;
      mem[464] = 16'b0000000000000000;
      mem[465] = 16'b0000000000000000;
      mem[466] = 16'b0000000000000000;
      mem[467] = 16'b0000000000000000;
      mem[468] = 16'b0000000000000000;
      mem[469] = 16'b0000000000000000;
      mem[470] = 16'b0000000000000000;
      mem[471] = 16'b0000000000000000;
      mem[472] = 16'b0000000000000000;
      mem[473] = 16'b0000000000000000;
      mem[474] = 16'b0000000000000000;
      mem[475] = 16'b0000000000000000;
      mem[476] = 16'b0000000000000000;
      mem[477] = 16'b0000000000000000;
      mem[478] = 16'b0000000000000000;
      mem[479] = 16'b0000000000000000;
      mem[480] = 16'b0000000000000000;
      mem[481] = 16'b0000000000000000;
      mem[482] = 16'b0000000000000000;
      mem[483] = 16'b0000000000000000;
      mem[484] = 16'b0000000000000000;
      mem[485] = 16'b0000000000000000;
      mem[486] = 16'b0000000000000000;
      mem[487] = 16'b0000000000000000;
      mem[488] = 16'b0000000000000000;
      mem[489] = 16'b0000000000000000;
      mem[490] = 16'b0000000000000000;
      mem[491] = 16'b0000000000000000;
      mem[492] = 16'b0000000000000000;
      mem[493] = 16'b0000000000000000;
      mem[494] = 16'b0000000000000000;
      mem[495] = 16'b0000000000000000;
      mem[496] = 16'b0000000000000000;
      mem[497] = 16'b0000000000000000;
      mem[498] = 16'b0000000000000000;
      mem[499] = 16'b0000000000000000;
      mem[500] = 16'b0000000000000000;
      mem[501] = 16'b0000000000000000;
      mem[502] = 16'b0000000000000000;
      mem[503] = 16'b0000000000000000;
      mem[504] = 16'b0000000000000000;
      mem[505] = 16'b0000000000000000;
      mem[506] = 16'b0000000000000000;
      mem[507] = 16'b0000000000000000;
      mem[508] = 16'b0000000000000000;
      mem[509] = 16'b0000000000000000;
      mem[510] = 16'b0000000000000000;
      mem[511] = 16'b0000000000000000;
      mem[512] = 16'b0000000000000000;
      mem[513] = 16'b0000000000000000;
      mem[514] = 16'b0000000000000000;
      mem[515] = 16'b0000000000000000;
      mem[516] = 16'b0000000000000000;
      mem[517] = 16'b0000000000000000;
      mem[518] = 16'b0000000000000000;
      mem[519] = 16'b0000000000000000;
      mem[520] = 16'b0000000000000000;
      mem[521] = 16'b0000000000000000;
      mem[522] = 16'b0000000000000000;
      mem[523] = 16'b0000000000000000;
      mem[524] = 16'b0000000000000000;
      mem[525] = 16'b0000000000000000;
      mem[526] = 16'b0000000000000000;
      mem[527] = 16'b0000000000000000;
      mem[528] = 16'b0000000000000000;
      mem[529] = 16'b0000000000000000;
      mem[530] = 16'b0000000000000000;
      mem[531] = 16'b0000000000000000;
      mem[532] = 16'b0000000000000000;
      mem[533] = 16'b0000000000000000;
      mem[534] = 16'b0000000000000000;
      mem[535] = 16'b0000000000000000;
      mem[536] = 16'b0000000000000000;
      mem[537] = 16'b0000000000000000;
      mem[538] = 16'b0000000000000000;
      mem[539] = 16'b0000000000000000;
      mem[540] = 16'b0000000000000000;
      mem[541] = 16'b0000000000000000;
      mem[542] = 16'b0000000000000000;
      mem[543] = 16'b0000000000000000;
      mem[544] = 16'b0000000000000000;
      mem[545] = 16'b0000000000000000;
      mem[546] = 16'b0000000000000000;
      mem[547] = 16'b0000000000000000;
      mem[548] = 16'b0000000000000000;
      mem[549] = 16'b0000000000000000;
      mem[550] = 16'b0000000000000000;
      mem[551] = 16'b0000000000000000;
      mem[552] = 16'b0000000000000000;
      mem[553] = 16'b0000000000000000;
      mem[554] = 16'b0000000000000000;
      mem[555] = 16'b0000000000000000;
      mem[556] = 16'b0000000000000000;
      mem[557] = 16'b0000000000000000;
      mem[558] = 16'b0000000000000000;
      mem[559] = 16'b0000000000000000;
      mem[560] = 16'b0000000000000000;
      mem[561] = 16'b0000000000000000;
      mem[562] = 16'b0000000000000000;
      mem[563] = 16'b0000000000000000;
      mem[564] = 16'b0000000000000000;
      mem[565] = 16'b0000000000000000;
      mem[566] = 16'b0000000000000000;
      mem[567] = 16'b0000000000000000;
      mem[568] = 16'b0000000000000000;
      mem[569] = 16'b0000000000000000;
      mem[570] = 16'b0000000000000000;
      mem[571] = 16'b0000000000000000;
      mem[572] = 16'b0000000000000000;
      mem[573] = 16'b0000000000000000;
      mem[574] = 16'b0000000000000000;
      mem[575] = 16'b0000000000000000;
      mem[576] = 16'b0000000000000000;
      mem[577] = 16'b0000000000000000;
      mem[578] = 16'b0000000000000000;
      mem[579] = 16'b0000000000000000;
      mem[580] = 16'b0000000000000000;
      mem[581] = 16'b0000000000000000;
      mem[582] = 16'b0000000000000000;
      mem[583] = 16'b0000000000000000;
      mem[584] = 16'b0000000000000000;
      mem[585] = 16'b0000000000000000;
      mem[586] = 16'b0000000000000000;
      mem[587] = 16'b0000000000000000;
      mem[588] = 16'b0000000000000000;
      mem[589] = 16'b0000000000000000;
      mem[590] = 16'b0000000000000000;
      mem[591] = 16'b0000000000000000;
      mem[592] = 16'b0000000000000000;
      mem[593] = 16'b0000000000000000;
      mem[594] = 16'b0000000000000000;
      mem[595] = 16'b0000000000000000;
      mem[596] = 16'b0000000000000000;
      mem[597] = 16'b0000000000000000;
      mem[598] = 16'b0000000000000000;
      mem[599] = 16'b0000000000000000;
      mem[600] = 16'b0000000000000000;
      mem[601] = 16'b0000000000000000;
      mem[602] = 16'b0000000000000000;
      mem[603] = 16'b0000000000000000;
      mem[604] = 16'b0000000000000000;
      mem[605] = 16'b0000000000000000;
      mem[606] = 16'b0000000000000000;
      mem[607] = 16'b0000000000000000;
      mem[608] = 16'b0000000000000000;
      mem[609] = 16'b0000000000000000;
      mem[610] = 16'b0000000000000000;
      mem[611] = 16'b0000000000000000;
      mem[612] = 16'b0000000000000000;
      mem[613] = 16'b0000000000000000;
      mem[614] = 16'b0000000000000000;
      mem[615] = 16'b0000000000000000;
      mem[616] = 16'b0000000000000000;
      mem[617] = 16'b0000000000000000;
      mem[618] = 16'b0000000000000000;
      mem[619] = 16'b0000000000000000;
      mem[620] = 16'b0000000000000000;
      mem[621] = 16'b0000000000000000;
      mem[622] = 16'b0000000000000000;
      mem[623] = 16'b0000000000000000;
      mem[624] = 16'b0000000000000000;
      mem[625] = 16'b0000000000000000;
      mem[626] = 16'b0000000000000000;
      mem[627] = 16'b0000000000000000;
      mem[628] = 16'b0000000000000000;
      mem[629] = 16'b0000000000000000;
      mem[630] = 16'b0000000000000000;
      mem[631] = 16'b0000000000000000;
      mem[632] = 16'b0000000000000000;
      mem[633] = 16'b0000000000000000;
      mem[634] = 16'b0000000000000000;
      mem[635] = 16'b0000000000000000;
      mem[636] = 16'b0000000000000000;
      mem[637] = 16'b0000000000000000;
      mem[638] = 16'b0000000000000000;
      mem[639] = 16'b0000000000000000;
      mem[640] = 16'b0000000000000000;
      mem[641] = 16'b0000000000000000;
      mem[642] = 16'b0000000000000000;
      mem[643] = 16'b0000000000000000;
      mem[644] = 16'b0000000000000000;
      mem[645] = 16'b0000000000000000;
      mem[646] = 16'b0000000000000000;
      mem[647] = 16'b0000000000000000;
      mem[648] = 16'b0000000000000000;
      mem[649] = 16'b0000000000000000;
      mem[650] = 16'b0000000000000000;
      mem[651] = 16'b0000000000000000;
      mem[652] = 16'b0000000000000000;
      mem[653] = 16'b0000000000000000;
      mem[654] = 16'b0000000000000000;
      mem[655] = 16'b0000000000000000;
      mem[656] = 16'b0000000000000000;
      mem[657] = 16'b0000000000000000;
      mem[658] = 16'b0000000000000000;
      mem[659] = 16'b0000000000000000;
      mem[660] = 16'b0000000000000000;
      mem[661] = 16'b0000000000000000;
      mem[662] = 16'b0000000000000000;
      mem[663] = 16'b0000000000000000;
      mem[664] = 16'b0000000000000000;
      mem[665] = 16'b0000000000000000;
      mem[666] = 16'b0000000000000000;
      mem[667] = 16'b0000000000000000;
      mem[668] = 16'b0000000000000000;
      mem[669] = 16'b0000000000000000;
      mem[670] = 16'b0000000000000000;
      mem[671] = 16'b0000000000000000;
      mem[672] = 16'b0000000000000000;
      mem[673] = 16'b0000000000000000;
      mem[674] = 16'b0000000000000000;
      mem[675] = 16'b0000000000000000;
      mem[676] = 16'b0000000000000000;
      mem[677] = 16'b0000000000000000;
      mem[678] = 16'b0000000000000000;
      mem[679] = 16'b0000000000000000;
      mem[680] = 16'b0000000000000000;
      mem[681] = 16'b0000000000000000;
      mem[682] = 16'b0000000000000000;
      mem[683] = 16'b0000000000000000;
      mem[684] = 16'b0000000000000000;
      mem[685] = 16'b0000000000000000;
      mem[686] = 16'b0000000000000000;
      mem[687] = 16'b0000000000000000;
      mem[688] = 16'b0000000000000000;
      mem[689] = 16'b0000000000000000;
      mem[690] = 16'b0000000000000000;
      mem[691] = 16'b0000000000000000;
      mem[692] = 16'b0000000000000000;
      mem[693] = 16'b0000000000000000;
      mem[694] = 16'b0000000000000000;
      mem[695] = 16'b0000000000000000;
      mem[696] = 16'b0000000000000000;
      mem[697] = 16'b0000000000000000;
      mem[698] = 16'b0000000000000000;
      mem[699] = 16'b0000000000000000;
      mem[700] = 16'b0000000000000000;
      mem[701] = 16'b0000000000000000;
      mem[702] = 16'b0000000000000000;
      mem[703] = 16'b0000000000000000;
      mem[704] = 16'b0000000000000000;
      mem[705] = 16'b0000000000000000;
      mem[706] = 16'b0000000000000000;
      mem[707] = 16'b0000000000000000;
      mem[708] = 16'b0000000000000000;
      mem[709] = 16'b0000000000000000;
      mem[710] = 16'b0000000000000000;
      mem[711] = 16'b0000000000000000;
      mem[712] = 16'b0000000000000000;
      mem[713] = 16'b0000000000000000;
      mem[714] = 16'b0000000000000000;
      mem[715] = 16'b0000000000000000;
      mem[716] = 16'b0000000000000000;
      mem[717] = 16'b0000000000000000;
      mem[718] = 16'b0000000000000000;
      mem[719] = 16'b0000000000000000;
      mem[720] = 16'b0000000000000000;
      mem[721] = 16'b0000000000000000;
      mem[722] = 16'b0000000000000000;
      mem[723] = 16'b0000000000000000;
      mem[724] = 16'b0000000000000000;
      mem[725] = 16'b0000000000000000;
      mem[726] = 16'b0000000000000000;
      mem[727] = 16'b0000000000000000;
      mem[728] = 16'b0000000000000000;
      mem[729] = 16'b0000000000000000;
      mem[730] = 16'b0000000000000000;
      mem[731] = 16'b0000000000000000;
      mem[732] = 16'b0000000000000000;
      mem[733] = 16'b0000000000000000;
      mem[734] = 16'b0000000000000000;
      mem[735] = 16'b0000000000000000;
      mem[736] = 16'b0000000000000000;
      mem[737] = 16'b0000000000000000;
      mem[738] = 16'b0000000000000000;
      mem[739] = 16'b0000000000000000;
      mem[740] = 16'b0000000000000000;
      mem[741] = 16'b0000000000000000;
      mem[742] = 16'b0000000000000000;
      mem[743] = 16'b0000000000000000;
      mem[744] = 16'b0000000000000000;
      mem[745] = 16'b0000000000000000;
      mem[746] = 16'b0000000000000000;
      mem[747] = 16'b0000000000000000;
      mem[748] = 16'b0000000000000000;
      mem[749] = 16'b0000000000000000;
      mem[750] = 16'b0000000000000000;
      mem[751] = 16'b0000000000000000;
      mem[752] = 16'b0000000000000000;
      mem[753] = 16'b0000000000000000;
      mem[754] = 16'b0000000000000000;
      mem[755] = 16'b0000000000000000;
      mem[756] = 16'b0000000000000000;
      mem[757] = 16'b0000000000000000;
      mem[758] = 16'b0000000000000000;
      mem[759] = 16'b0000000000000000;
      mem[760] = 16'b0000000000000000;
      mem[761] = 16'b0000000000000000;
      mem[762] = 16'b0000000000000000;
      mem[763] = 16'b0000000000000000;
      mem[764] = 16'b0000000000000000;
      mem[765] = 16'b0000000000000000;
      mem[766] = 16'b0000000000000000;
      mem[767] = 16'b0000000000000000;
      mem[768] = 16'b0000000000000000;
      mem[769] = 16'b0000000000000000;
      mem[770] = 16'b0000000000000000;
      mem[771] = 16'b0000000000000000;
      mem[772] = 16'b0000000000000000;
      mem[773] = 16'b0000000000000000;
      mem[774] = 16'b0000000000000000;
      mem[775] = 16'b0000000000000000;
      mem[776] = 16'b0000000000000000;
      mem[777] = 16'b0000000000000000;
      mem[778] = 16'b0000000000000000;
      mem[779] = 16'b0000000000000000;
      mem[780] = 16'b0000000000000000;
      mem[781] = 16'b0000000000000000;
      mem[782] = 16'b0000000000000000;
      mem[783] = 16'b0000000000000000;
      mem[784] = 16'b0000000000000000;
      mem[785] = 16'b0000000000000000;
      mem[786] = 16'b0000000000000000;
      mem[787] = 16'b0000000000000000;
      mem[788] = 16'b0000000000000000;
      mem[789] = 16'b0000000000000000;
      mem[790] = 16'b0000000000000000;
      mem[791] = 16'b0000000000000000;
      mem[792] = 16'b0000000000000000;
      mem[793] = 16'b0000000000000000;
      mem[794] = 16'b0000000000000000;
      mem[795] = 16'b0000000000000000;
      mem[796] = 16'b0000000000000000;
      mem[797] = 16'b0000000000000000;
      mem[798] = 16'b0000000000000000;
      mem[799] = 16'b0000000000000000;
      mem[800] = 16'b0000000000000000;
      mem[801] = 16'b0000000000000000;
      mem[802] = 16'b0000000000000000;
      mem[803] = 16'b0000000000000000;
      mem[804] = 16'b0000000000000000;
      mem[805] = 16'b0000000000000000;
      mem[806] = 16'b0000000000000000;
      mem[807] = 16'b0000000000000000;
      mem[808] = 16'b0000000000000000;
      mem[809] = 16'b0000000000000000;
      mem[810] = 16'b0000000000000000;
      mem[811] = 16'b0000000000000000;
      mem[812] = 16'b0000000000000000;
      mem[813] = 16'b0000000000000000;
      mem[814] = 16'b0000000000000000;
      mem[815] = 16'b0000000000000000;
      mem[816] = 16'b0000000000000000;
      mem[817] = 16'b0000000000000000;
      mem[818] = 16'b0000000000000000;
      mem[819] = 16'b0000000000000000;
      mem[820] = 16'b0000000000000000;
      mem[821] = 16'b0000000000000000;
      mem[822] = 16'b0000000000000000;
      mem[823] = 16'b0000000000000000;
      mem[824] = 16'b0000000000000000;
      mem[825] = 16'b0000000000000000;
      mem[826] = 16'b0000000000000000;
      mem[827] = 16'b0000000000000000;
      mem[828] = 16'b0000000000000000;
      mem[829] = 16'b0000000000000000;
      mem[830] = 16'b0000000000000000;
      mem[831] = 16'b0000000000000000;
      mem[832] = 16'b0000000000000000;
      mem[833] = 16'b0000000000000000;
      mem[834] = 16'b0000000000000000;
      mem[835] = 16'b0000000000000000;
      mem[836] = 16'b0000000000000000;
      mem[837] = 16'b0000000000000000;
      mem[838] = 16'b0000000000000000;
      mem[839] = 16'b0000000000000000;
      mem[840] = 16'b0000000000000000;
      mem[841] = 16'b0000000000000000;
      mem[842] = 16'b0000000000000000;
      mem[843] = 16'b0000000000000000;
      mem[844] = 16'b0000000000000000;
      mem[845] = 16'b0000000000000000;
      mem[846] = 16'b0000000000000000;
      mem[847] = 16'b0000000000000000;
      mem[848] = 16'b0000000000000000;
      mem[849] = 16'b0000000000000000;
      mem[850] = 16'b0000000000000000;
      mem[851] = 16'b0000000000000000;
      mem[852] = 16'b0000000000000000;
      mem[853] = 16'b0000000000000000;
      mem[854] = 16'b0000000000000000;
      mem[855] = 16'b0000000000000000;
      mem[856] = 16'b0000000000000000;
      mem[857] = 16'b0000000000000000;
      mem[858] = 16'b0000000000000000;
      mem[859] = 16'b0000000000000000;
      mem[860] = 16'b0000000000000000;
      mem[861] = 16'b0000000000000000;
      mem[862] = 16'b0000000000000000;
      mem[863] = 16'b0000000000000000;
      mem[864] = 16'b0000000000000000;
      mem[865] = 16'b0000000000000000;
      mem[866] = 16'b0000000000000000;
      mem[867] = 16'b0000000000000000;
      mem[868] = 16'b0000000000000000;
      mem[869] = 16'b0000000000000000;
      mem[870] = 16'b0000000000000000;
      mem[871] = 16'b0000000000000000;
      mem[872] = 16'b0000000000000000;
      mem[873] = 16'b0000000000000000;
      mem[874] = 16'b0000000000000000;
      mem[875] = 16'b0000000000000000;
      mem[876] = 16'b0000000000000000;
      mem[877] = 16'b0000000000000000;
      mem[878] = 16'b0000000000000000;
      mem[879] = 16'b0000000000000000;
      mem[880] = 16'b0000000000000000;
      mem[881] = 16'b0000000000000000;
      mem[882] = 16'b0000000000000000;
      mem[883] = 16'b0000000000000000;
      mem[884] = 16'b0000000000000000;
      mem[885] = 16'b0000000000000000;
      mem[886] = 16'b0000000000000000;
      mem[887] = 16'b0000000000000000;
      mem[888] = 16'b0000000000000000;
      mem[889] = 16'b0000000000000000;
      mem[890] = 16'b0000000000000000;
      mem[891] = 16'b0000000000000000;
      mem[892] = 16'b0000000000000000;
      mem[893] = 16'b0000000000000000;
      mem[894] = 16'b0000000000000000;
      mem[895] = 16'b0000000000000000;
      mem[896] = 16'b0000000000000000;
      mem[897] = 16'b0000000000000000;
      mem[898] = 16'b0000000000000000;
      mem[899] = 16'b0000000000000000;
      mem[900] = 16'b0000000000000000;
      mem[901] = 16'b0000000000000000;
      mem[902] = 16'b0000000000000000;
      mem[903] = 16'b0000000000000000;
      mem[904] = 16'b0000000000000000;
      mem[905] = 16'b0000000000000000;
      mem[906] = 16'b0000000000000000;
      mem[907] = 16'b0000000000000000;
      mem[908] = 16'b0000000000000000;
      mem[909] = 16'b0000000000000000;
      mem[910] = 16'b0000000000000000;
      mem[911] = 16'b0000000000000000;
      mem[912] = 16'b0000000000000000;
      mem[913] = 16'b0000000000000000;
      mem[914] = 16'b0000000000000000;
      mem[915] = 16'b0000000000000000;
      mem[916] = 16'b0000000000000000;
      mem[917] = 16'b0000000000000000;
      mem[918] = 16'b0000000000000000;
      mem[919] = 16'b0000000000000000;
      mem[920] = 16'b0000000000000000;
      mem[921] = 16'b0000000000000000;
      mem[922] = 16'b0000000000000000;
      mem[923] = 16'b0000000000000000;
      mem[924] = 16'b0000000000000000;
      mem[925] = 16'b0000000000000000;
      mem[926] = 16'b0000000000000000;
      mem[927] = 16'b0000000000000000;
      mem[928] = 16'b0000000000000000;
      mem[929] = 16'b0000000000000000;
      mem[930] = 16'b0000000000000000;
      mem[931] = 16'b0000000000000000;
      mem[932] = 16'b0000000000000000;
      mem[933] = 16'b0000000000000000;
      mem[934] = 16'b0000000000000000;
      mem[935] = 16'b0000000000000000;
      mem[936] = 16'b0000000000000000;
      mem[937] = 16'b0000000000000000;
      mem[938] = 16'b0000000000000000;
      mem[939] = 16'b0000000000000000;
      mem[940] = 16'b0000000000000000;
      mem[941] = 16'b0000000000000000;
      mem[942] = 16'b0000000000000000;
      mem[943] = 16'b0000000000000000;
      mem[944] = 16'b0000000000000000;
      mem[945] = 16'b0000000000000000;
      mem[946] = 16'b0000000000000000;
      mem[947] = 16'b0000000000000000;
      mem[948] = 16'b0000000000000000;
      mem[949] = 16'b0000000000000000;
      mem[950] = 16'b0000000000000000;
      mem[951] = 16'b0000000000000000;
      mem[952] = 16'b0000000000000000;
      mem[953] = 16'b0000000000000000;
      mem[954] = 16'b0000000000000000;
      mem[955] = 16'b0000000000000000;
      mem[956] = 16'b0000000000000000;
      mem[957] = 16'b0000000000000000;
      mem[958] = 16'b0000000000000000;
      mem[959] = 16'b0000000000000000;
      mem[960] = 16'b0000000000000000;
      mem[961] = 16'b0000000000000000;
      mem[962] = 16'b0000000000000000;
      mem[963] = 16'b0000000000000000;
      mem[964] = 16'b0000000000000000;
      mem[965] = 16'b0000000000000000;
      mem[966] = 16'b0000000000000000;
      mem[967] = 16'b0000000000000000;
      mem[968] = 16'b0000000000000000;
      mem[969] = 16'b0000000000000000;
      mem[970] = 16'b0000000000000000;
      mem[971] = 16'b0000000000000000;
      mem[972] = 16'b0000000000000000;
      mem[973] = 16'b0000000000000000;
      mem[974] = 16'b0000000000000000;
      mem[975] = 16'b0000000000000000;
      mem[976] = 16'b0000000000000000;
      mem[977] = 16'b0000000000000000;
      mem[978] = 16'b0000000000000000;
      mem[979] = 16'b0000000000000000;
      mem[980] = 16'b0000000000000000;
      mem[981] = 16'b0000000000000000;
      mem[982] = 16'b0000000000000000;
      mem[983] = 16'b0000000000000000;
      mem[984] = 16'b0000000000000000;
      mem[985] = 16'b0000000000000000;
      mem[986] = 16'b0000000000000000;
      mem[987] = 16'b0000000000000000;
      mem[988] = 16'b0000000000000000;
      mem[989] = 16'b0000000000000000;
      mem[990] = 16'b0000000000000000;
      mem[991] = 16'b0000000000000000;
      mem[992] = 16'b0000000000000000;
      mem[993] = 16'b0000000000000000;
      mem[994] = 16'b0000000000000000;
      mem[995] = 16'b0000000000000000;
      mem[996] = 16'b0000000000000000;
      mem[997] = 16'b0000000000000000;
      mem[998] = 16'b0000000000000000;
      mem[999] = 16'b0000000000000000;
      mem[1000] = 16'b0000000000000000;
      mem[1001] = 16'b0000000000000000;
      mem[1002] = 16'b0000000000000000;
      mem[1003] = 16'b0000000000000000;
      mem[1004] = 16'b0000000000000000;
      mem[1005] = 16'b0000000000000000;
      mem[1006] = 16'b0000000000000000;
      mem[1007] = 16'b0000000000000000;
      mem[1008] = 16'b0000000000000000;
      mem[1009] = 16'b0000000000000000;
      mem[1010] = 16'b0000000000000000;
      mem[1011] = 16'b0000000000000000;
      mem[1012] = 16'b0000000000000000;
      mem[1013] = 16'b0000000000000000;
      mem[1014] = 16'b0000000000000000;
      mem[1015] = 16'b0000000000000000;
      mem[1016] = 16'b0000000000000000;
      mem[1017] = 16'b0000000000000000;
      mem[1018] = 16'b0000000000000000;
      mem[1019] = 16'b0000000000000000;
      mem[1020] = 16'b0000000000000000;
      mem[1021] = 16'b0000000000000000;
      mem[1022] = 16'b0000000000000000;
      mem[1023] = 16'b0000000000000000;
   end
   assign read_addr = i[9:0];
   assign write_addr = i[19:10];
   assign write_value = i[35:20];
   assign write_enable = i[36:36];
   assign clock = clock_reset[0:0];
   always @(posedge clock) begin
      o <= mem[read_addr];
   end
   always @(posedge clock) begin
      if (write_enable) begin
         mem[write_addr] <= write_value;
      end
   end
endmodule
module top_T1(input wire [1:0] clock_reset, input wire [17:0] i, output wire [31:0] o);
   wire [47:0] od;
   wire [15:0] d;
   wire [15:0] q;
   assign o = od[31:0];
   top_T1_memory c0(.clock_reset(clock_reset), .i(d[15:0]), .o(q[15:0]));
   assign d = od[47:32];
   assign od = kernel_reg_ker(clock_reset, i, q);
   function [47:0] kernel_reg_ker(input reg [1:0] arg_0, input reg [17:0] arg_1, input reg [15:0] arg_2);
         reg [0:0] or0;
         reg [17:0] or1;
         reg [0:0] or2;
         reg [0:0] or3;
         reg [0:0] or4;
         reg [15:0] or5;
         reg [15:0] or6;
         reg [0:0] or7;
         reg [15:0] or8;
         reg [31:0] or9;
         reg [0:0] or10;
         reg [15:0] or11;
         reg [15:0] or12;
         reg [15:0] or13;
         reg [47:0] or14;
         reg [1:0] or15;
         localparam ol0 = 16'b0000000000000000;
         localparam ol1 = 16'b0000000000000000;
         localparam ol2 = 16'b0000000000000000;
         begin
            or15 = arg_0;
            or1 = arg_1;
            or5 = arg_2;
            or0 = or1[16:16];
            or2 = or1[17:17];
            or3 = ~or2;
            or4 = or0 & or3;
            or6 = or4 ? or5 : ol0;
            or7 = or1[16:16];
            or8 = or7 ? or5 : ol1;
            or9 = {or8, or6};
            or10 = or1[17:17];
            or11 = or1[15:0];
            or12 = or10 ? or11 : or5;
            or13 = ol2;
            or13[15:0] = or12;
            or14 = {or13, or9};
            kernel_reg_ker = or14;
         end
   endfunction
endmodule
module top_T1_memory(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000101;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000101;
      end else begin
         o <= i;
      end
   end
endmodule
module top_T2(input wire [1:0] clock_reset, input wire [17:0] i, output wire [31:0] o);
   wire [47:0] od;
   wire [15:0] d;
   wire [15:0] q;
   assign o = od[31:0];
   top_T2_memory c0(.clock_reset(clock_reset), .i(d[15:0]), .o(q[15:0]));
   assign d = od[47:32];
   assign od = kernel_reg_ker(clock_reset, i, q);
   function [47:0] kernel_reg_ker(input reg [1:0] arg_0, input reg [17:0] arg_1, input reg [15:0] arg_2);
         reg [0:0] or0;
         reg [17:0] or1;
         reg [0:0] or2;
         reg [0:0] or3;
         reg [0:0] or4;
         reg [15:0] or5;
         reg [15:0] or6;
         reg [0:0] or7;
         reg [15:0] or8;
         reg [31:0] or9;
         reg [0:0] or10;
         reg [15:0] or11;
         reg [15:0] or12;
         reg [15:0] or13;
         reg [47:0] or14;
         reg [1:0] or15;
         localparam ol0 = 16'b0000000000000000;
         localparam ol1 = 16'b0000000000000000;
         localparam ol2 = 16'b0000000000000000;
         begin
            or15 = arg_0;
            or1 = arg_1;
            or5 = arg_2;
            or0 = or1[16:16];
            or2 = or1[17:17];
            or3 = ~or2;
            or4 = or0 & or3;
            or6 = or4 ? or5 : ol0;
            or7 = or1[16:16];
            or8 = or7 ? or5 : ol1;
            or9 = {or8, or6};
            or10 = or1[17:17];
            or11 = or1[15:0];
            or12 = or10 ? or11 : or5;
            or13 = ol2;
            or13[15:0] = or12;
            or14 = {or13, or9};
            kernel_reg_ker = or14;
         end
   endfunction
endmodule
module top_T2_memory(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_regs(input wire [1:0] clock_reset, input wire [20:0] i, output wire [15:0] o);
   wire [143:0] od;
   wire [127:0] d;
   wire [127:0] q;
   assign o = od[15:0];
   top_regs_rg c0(.clock_reset(clock_reset), .i(d[127:0]), .o(q[127:0]));
   assign d = od[143:16];
   assign od = kernel_reg_file(clock_reset, i, q);
   function [143:0] kernel_reg_file(input reg [1:0] arg_0, input reg [20:0] arg_1, input reg [127:0] arg_2);
         reg [127:0] or0;
         // d
         reg [127:0] or1;
         reg [17:0] or2;
         reg [20:0] or3;
         reg [0:0] or4;
         reg [17:0] or5;
         reg [0:0] or6;
         reg [0:0] or7;
         reg [0:0] or8;
         reg [2:0] or9;
         reg [15:0] or10;
         reg [15:0] or11;
         reg [15:0] or12;
         reg [15:0] or13;
         reg [15:0] or14;
         reg [15:0] or15;
         reg [15:0] or16;
         reg [15:0] or17;
         reg [15:0] or18;
         reg [15:0] or19;
         reg [17:0] or20;
         reg [0:0] or21;
         reg [2:0] or22;
         reg [17:0] or23;
         reg [15:0] or24;
         // d
         reg [127:0] or25;
         reg [17:0] or26;
         reg [15:0] or27;
         // d
         reg [127:0] or28;
         reg [17:0] or29;
         reg [15:0] or30;
         // d
         reg [127:0] or31;
         reg [17:0] or32;
         reg [15:0] or33;
         // d
         reg [127:0] or34;
         reg [17:0] or35;
         reg [15:0] or36;
         // d
         reg [127:0] or37;
         reg [17:0] or38;
         reg [15:0] or39;
         // d
         reg [127:0] or40;
         reg [17:0] or41;
         reg [15:0] or42;
         // d
         reg [127:0] or43;
         reg [17:0] or44;
         reg [15:0] or45;
         // d
         reg [127:0] or46;
         // d
         reg [127:0] or47;
         // d
         reg [127:0] or48;
         reg [143:0] or49;
         reg [1:0] or50;
         localparam ol0 = 128'bXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX;
         localparam ol1 = 3'b000;
         localparam ol2 = 3'b001;
         localparam ol3 = 3'b010;
         localparam ol4 = 3'b011;
         localparam ol5 = 3'b100;
         localparam ol6 = 3'b101;
         localparam ol7 = 3'b110;
         localparam ol8 = 3'b111;
         localparam ol9 = 16'b0000000000000000;
         localparam ol10 = 3'b000;
         localparam ol11 = 3'b001;
         localparam ol12 = 3'b010;
         localparam ol13 = 3'b011;
         localparam ol14 = 3'b100;
         localparam ol15 = 3'b101;
         localparam ol16 = 3'b110;
         localparam ol17 = 3'b111;
         begin
            or50 = arg_0;
            or3 = arg_1;
            or0 = arg_2;
            or1 = ol0;
            or1[127:0] = or0;
            or2 = or3[17:0];
            or4 = or2[16:16];
            or5 = or3[17:0];
            or6 = or5[17:17];
            or7 = ~or6;
            or8 = or4 & or7;
            or9 = or3[20:18];
            or10 = or0[15:0];
            or11 = or0[31:16];
            or12 = or0[47:32];
            or13 = or0[63:48];
            or14 = or0[79:64];
            or15 = or0[95:80];
            or16 = or0[111:96];
            or17 = or0[127:112];
            case (or9)
               3'b000 : or18 = or10;
               3'b001 : or18 = or11;
               3'b010 : or18 = or12;
               3'b011 : or18 = or13;
               3'b100 : or18 = or14;
               3'b101 : or18 = or15;
               3'b110 : or18 = or16;
               3'b111 : or18 = or17;
            endcase
            or19 = or8 ? or18 : ol9;
            or20 = or3[17:0];
            or21 = or20[17:17];
            or22 = or3[20:18];
            or23 = or3[17:0];
            or24 = or23[15:0];
            or25 = or1;
            or25[15:0] = or24;
            or26 = or3[17:0];
            or27 = or26[15:0];
            or28 = or1;
            or28[31:16] = or27;
            or29 = or3[17:0];
            or30 = or29[15:0];
            or31 = or1;
            or31[47:32] = or30;
            or32 = or3[17:0];
            or33 = or32[15:0];
            or34 = or1;
            or34[63:48] = or33;
            or35 = or3[17:0];
            or36 = or35[15:0];
            or37 = or1;
            or37[79:64] = or36;
            or38 = or3[17:0];
            or39 = or38[15:0];
            or40 = or1;
            or40[95:80] = or39;
            or41 = or3[17:0];
            or42 = or41[15:0];
            or43 = or1;
            or43[111:96] = or42;
            or44 = or3[17:0];
            or45 = or44[15:0];
            or46 = or1;
            or46[127:112] = or45;
            case (or22)
               3'b000 : or47 = or25;
               3'b001 : or47 = or28;
               3'b010 : or47 = or31;
               3'b011 : or47 = or34;
               3'b100 : or47 = or37;
               3'b101 : or47 = or40;
               3'b110 : or47 = or43;
               3'b111 : or47 = or46;
            endcase
            or48 = or21 ? or47 : or1;
            or49 = {or48, or19};
            kernel_reg_file = or49;
         end
   endfunction
endmodule
module top_regs_rg(input wire [1:0] clock_reset, input wire [127:0] i, output wire [127:0] o);
   top_regs_rg_0 c0(.clock_reset(clock_reset), .i(i[15:0]), .o(o[15:0]));
   top_regs_rg_1 c1(.clock_reset(clock_reset), .i(i[31:16]), .o(o[31:16]));
   top_regs_rg_2 c2(.clock_reset(clock_reset), .i(i[47:32]), .o(o[47:32]));
   top_regs_rg_3 c3(.clock_reset(clock_reset), .i(i[63:48]), .o(o[63:48]));
   top_regs_rg_4 c4(.clock_reset(clock_reset), .i(i[79:64]), .o(o[79:64]));
   top_regs_rg_5 c5(.clock_reset(clock_reset), .i(i[95:80]), .o(o[95:80]));
   top_regs_rg_6 c6(.clock_reset(clock_reset), .i(i[111:96]), .o(o[111:96]));
   top_regs_rg_7 c7(.clock_reset(clock_reset), .i(i[127:112]), .o(o[127:112]));
endmodule
module top_regs_rg_0(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_regs_rg_1(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_regs_rg_2(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_regs_rg_3(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_regs_rg_4(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_regs_rg_5(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_regs_rg_6(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
module top_regs_rg_7(input wire [1:0] clock_reset, input wire [15:0] i, output reg [15:0] o);
   wire  clock;
   wire  reset;
   assign clock = clock_reset[0];
   assign reset = clock_reset[1];
   initial begin
      o = 16'b0000000000000000;
   end
   always @(posedge clock) begin
      if (reset) begin
         o <= 16'b0000000000000000;
      end else begin
         o <= i;
      end
   end
endmodule
