module top(input wire [1:0] clock_reset, input wire [7:0] i, output wire [4:0] o);
   assign o = kernel_adder_4bit(clock_reset, i);
   function [4:0] kernel_adder_4bit(input reg [1:0] arg_0, input reg [7:0] arg_1);
         reg [3:0] or0;
         reg [7:0] or1;
         reg [0:0] or2;
         reg [3:0] or3;
         reg [0:0] or4;
         reg [2:0] or5;
         reg [2:0] or6;
         reg [2:0] or7;
         reg [0:0] or8;
         reg [0:0] or9;
         reg [1:0] or10;
         reg [1:0] or11;
         reg [0:0] or12;
         reg [0:0] or13;
         reg [1:0] or14;
         reg [0:0] or15;
         reg [0:0] or16;
         reg [0:0] or17;
         reg [0:0] or18;
         reg [0:0] or19;
         reg [1:0] or20;
         reg [0:0] or21;
         reg [0:0] or22;
         reg [0:0] or23;
         reg [1:0] or24;
         reg [1:0] or25;
         reg [0:0] or26;
         reg [0:0] or27;
         reg [0:0] or28;
         reg [1:0] or29;
         reg [1:0] or30;
         reg [0:0] or31;
         reg [0:0] or32;
         reg [1:0] or33;
         reg [0:0] or34;
         reg [0:0] or35;
         reg [0:0] or36;
         reg [0:0] or37;
         reg [0:0] or38;
         reg [1:0] or39;
         reg [0:0] or40;
         reg [0:0] or41;
         reg [0:0] or42;
         reg [1:0] or43;
         reg [1:0] or44;
         reg [0:0] or45;
         reg [0:0] or46;
         reg [1:0] or47;
         reg [0:0] or48;
         reg [0:0] or49;
         reg [0:0] or50;
         reg [1:0] or51;
         reg [1:0] or52;
         reg [1:0] or53;
         reg [0:0] or54;
         reg [0:0] or55;
         reg [3:0] or56;
         reg [0:0] or57;
         reg [3:0] or58;
         reg [0:0] or59;
         reg [2:0] or60;
         reg [2:0] or61;
         reg [2:0] or62;
         reg [0:0] or63;
         reg [0:0] or64;
         reg [1:0] or65;
         reg [1:0] or66;
         reg [0:0] or67;
         reg [0:0] or68;
         reg [1:0] or69;
         reg [0:0] or70;
         reg [0:0] or71;
         reg [0:0] or72;
         reg [0:0] or73;
         reg [0:0] or74;
         reg [1:0] or75;
         reg [0:0] or76;
         reg [0:0] or77;
         reg [0:0] or78;
         reg [1:0] or79;
         reg [1:0] or80;
         reg [0:0] or81;
         reg [0:0] or82;
         reg [0:0] or83;
         reg [1:0] or84;
         reg [1:0] or85;
         reg [0:0] or86;
         reg [0:0] or87;
         reg [1:0] or88;
         reg [0:0] or89;
         reg [0:0] or90;
         reg [0:0] or91;
         reg [0:0] or92;
         reg [0:0] or93;
         reg [1:0] or94;
         reg [0:0] or95;
         reg [0:0] or96;
         reg [0:0] or97;
         reg [1:0] or98;
         reg [1:0] or99;
         reg [0:0] or100;
         reg [0:0] or101;
         reg [1:0] or102;
         reg [0:0] or103;
         reg [0:0] or104;
         reg [0:0] or105;
         reg [1:0] or106;
         reg [1:0] or107;
         reg [0:0] or108;
         reg [0:0] or109;
         reg [3:0] or110;
         reg [0:0] or111;
         reg [3:0] or112;
         reg [0:0] or113;
         reg [2:0] or114;
         reg [2:0] or115;
         reg [2:0] or116;
         reg [0:0] or117;
         reg [0:0] or118;
         reg [1:0] or119;
         reg [1:0] or120;
         reg [0:0] or121;
         reg [0:0] or122;
         reg [1:0] or123;
         reg [0:0] or124;
         reg [0:0] or125;
         reg [0:0] or126;
         reg [0:0] or127;
         reg [0:0] or128;
         reg [1:0] or129;
         reg [0:0] or130;
         reg [0:0] or131;
         reg [0:0] or132;
         reg [1:0] or133;
         reg [1:0] or134;
         reg [0:0] or135;
         reg [0:0] or136;
         reg [0:0] or137;
         reg [1:0] or138;
         reg [1:0] or139;
         reg [0:0] or140;
         reg [0:0] or141;
         reg [1:0] or142;
         reg [0:0] or143;
         reg [0:0] or144;
         reg [0:0] or145;
         reg [0:0] or146;
         reg [0:0] or147;
         reg [1:0] or148;
         reg [0:0] or149;
         reg [0:0] or150;
         reg [0:0] or151;
         reg [1:0] or152;
         reg [1:0] or153;
         reg [0:0] or154;
         reg [0:0] or155;
         reg [1:0] or156;
         reg [0:0] or157;
         reg [0:0] or158;
         reg [0:0] or159;
         reg [1:0] or160;
         reg [1:0] or161;
         reg [0:0] or162;
         reg [0:0] or163;
         reg [3:0] or164;
         reg [0:0] or165;
         reg [3:0] or166;
         reg [0:0] or167;
         reg [2:0] or168;
         reg [2:0] or169;
         reg [2:0] or170;
         reg [0:0] or171;
         reg [0:0] or172;
         reg [1:0] or173;
         reg [1:0] or174;
         reg [0:0] or175;
         reg [0:0] or176;
         reg [1:0] or177;
         reg [0:0] or178;
         reg [0:0] or179;
         reg [0:0] or180;
         reg [0:0] or181;
         reg [0:0] or182;
         reg [1:0] or183;
         reg [0:0] or184;
         reg [0:0] or185;
         reg [0:0] or186;
         reg [1:0] or187;
         reg [1:0] or188;
         reg [0:0] or189;
         reg [0:0] or190;
         reg [0:0] or191;
         reg [1:0] or192;
         reg [1:0] or193;
         reg [0:0] or194;
         reg [0:0] or195;
         reg [1:0] or196;
         reg [0:0] or197;
         reg [0:0] or198;
         reg [0:0] or199;
         reg [0:0] or200;
         reg [0:0] or201;
         reg [1:0] or202;
         reg [0:0] or203;
         reg [0:0] or204;
         reg [0:0] or205;
         reg [1:0] or206;
         reg [1:0] or207;
         reg [0:0] or208;
         reg [0:0] or209;
         reg [1:0] or210;
         reg [0:0] or211;
         reg [0:0] or212;
         reg [0:0] or213;
         reg [1:0] or214;
         reg [1:0] or215;
         reg [0:0] or216;
         reg [0:0] or217;
         reg [4:0] or218;
         localparam ol0 = 3'b000;
         localparam ol1 = 1'b0;
         localparam ol2 = 2'b00;
         localparam ol3 = 2'b00;
         localparam ol4 = 2'b00;
         localparam ol5 = 2'b00;
         localparam ol6 = 2'b00;
         localparam ol7 = 3'b000;
         localparam ol8 = 2'b00;
         localparam ol9 = 2'b00;
         localparam ol10 = 2'b00;
         localparam ol11 = 2'b00;
         localparam ol12 = 2'b00;
         localparam ol13 = 3'b000;
         localparam ol14 = 2'b00;
         localparam ol15 = 2'b00;
         localparam ol16 = 2'b00;
         localparam ol17 = 2'b00;
         localparam ol18 = 2'b00;
         localparam ol19 = 3'b000;
         localparam ol20 = 2'b00;
         localparam ol21 = 2'b00;
         localparam ol22 = 2'b00;
         localparam ol23 = 2'b00;
         localparam ol24 = 2'b00;
         begin
            or53 = arg_0;
            or1 = arg_1;
            or0 = or1[3:0];
            or2 = or0[3:3];
            or3 = or1[7:4];
            or4 = or3[3:3];
            or5 = ol0;
            or5[0:0] = or2;
            or6 = or5;
            or6[1:1] = or4;
            or7 = or6;
            or7[2:2] = ol1;
            or8 = or7[0:0];
            or9 = or7[1:1];
            or10 = ol2;
            or10[0:0] = or8;
            or11 = or10;
            or11[1:1] = or9;
            or12 = or11[0:0];
            or13 = or11[1:1];
            or14 = {or13, or12};
            or15 = or14[0:0];
            or16 = or14[1:1];
            or17 = or15 ^ or16;
            or18 = or11[0:0];
            or19 = or11[1:1];
            or20 = {or19, or18};
            or21 = or20[0:0];
            or22 = or20[1:1];
            or23 = or21 & or22;
            or24 = ol3;
            or24[0:0] = or17;
            or25 = or24;
            or25[1:1] = or23;
            or26 = or25[0:0];
            or27 = or25[1:1];
            or28 = or7[2:2];
            or29 = ol4;
            or29[0:0] = or28;
            or30 = or29;
            or30[1:1] = or26;
            or31 = or30[0:0];
            or32 = or30[1:1];
            or33 = {or32, or31};
            or34 = or33[0:0];
            or35 = or33[1:1];
            or36 = or34 ^ or35;
            or37 = or30[0:0];
            or38 = or30[1:1];
            or39 = {or38, or37};
            or40 = or39[0:0];
            or41 = or39[1:1];
            or42 = or40 & or41;
            or43 = ol5;
            or43[0:0] = or36;
            or44 = or43;
            or44[1:1] = or42;
            or45 = or44[0:0];
            or46 = or44[1:1];
            or47 = {or46, or27};
            or48 = or47[1:1];
            or49 = or47[0:0];
            or50 = or48 | or49;
            or51 = ol6;
            or51[0:0] = or45;
            or52 = or51;
            or52[1:1] = or50;
            or54 = or52[0:0];
            or55 = or52[1:1];
            or56 = or1[3:0];
            or57 = or56[2:2];
            or58 = or1[7:4];
            or59 = or58[2:2];
            or60 = ol7;
            or60[0:0] = or57;
            or61 = or60;
            or61[1:1] = or59;
            or62 = or61;
            or62[2:2] = or55;
            or63 = or62[0:0];
            or64 = or62[1:1];
            or65 = ol8;
            or65[0:0] = or63;
            or66 = or65;
            or66[1:1] = or64;
            or67 = or66[0:0];
            or68 = or66[1:1];
            or69 = {or68, or67};
            or70 = or69[0:0];
            or71 = or69[1:1];
            or72 = or70 ^ or71;
            or73 = or66[0:0];
            or74 = or66[1:1];
            or75 = {or74, or73};
            or76 = or75[0:0];
            or77 = or75[1:1];
            or78 = or76 & or77;
            or79 = ol9;
            or79[0:0] = or72;
            or80 = or79;
            or80[1:1] = or78;
            or81 = or80[0:0];
            or82 = or80[1:1];
            or83 = or62[2:2];
            or84 = ol10;
            or84[0:0] = or83;
            or85 = or84;
            or85[1:1] = or81;
            or86 = or85[0:0];
            or87 = or85[1:1];
            or88 = {or87, or86};
            or89 = or88[0:0];
            or90 = or88[1:1];
            or91 = or89 ^ or90;
            or92 = or85[0:0];
            or93 = or85[1:1];
            or94 = {or93, or92};
            or95 = or94[0:0];
            or96 = or94[1:1];
            or97 = or95 & or96;
            or98 = ol11;
            or98[0:0] = or91;
            or99 = or98;
            or99[1:1] = or97;
            or100 = or99[0:0];
            or101 = or99[1:1];
            or102 = {or101, or82};
            or103 = or102[1:1];
            or104 = or102[0:0];
            or105 = or103 | or104;
            or106 = ol12;
            or106[0:0] = or100;
            or107 = or106;
            or107[1:1] = or105;
            or108 = or107[0:0];
            or109 = or107[1:1];
            or110 = or1[3:0];
            or111 = or110[1:1];
            or112 = or1[7:4];
            or113 = or112[1:1];
            or114 = ol13;
            or114[0:0] = or111;
            or115 = or114;
            or115[1:1] = or113;
            or116 = or115;
            or116[2:2] = or109;
            or117 = or116[0:0];
            or118 = or116[1:1];
            or119 = ol14;
            or119[0:0] = or117;
            or120 = or119;
            or120[1:1] = or118;
            or121 = or120[0:0];
            or122 = or120[1:1];
            or123 = {or122, or121};
            or124 = or123[0:0];
            or125 = or123[1:1];
            or126 = or124 ^ or125;
            or127 = or120[0:0];
            or128 = or120[1:1];
            or129 = {or128, or127};
            or130 = or129[0:0];
            or131 = or129[1:1];
            or132 = or130 & or131;
            or133 = ol15;
            or133[0:0] = or126;
            or134 = or133;
            or134[1:1] = or132;
            or135 = or134[0:0];
            or136 = or134[1:1];
            or137 = or116[2:2];
            or138 = ol16;
            or138[0:0] = or137;
            or139 = or138;
            or139[1:1] = or135;
            or140 = or139[0:0];
            or141 = or139[1:1];
            or142 = {or141, or140};
            or143 = or142[0:0];
            or144 = or142[1:1];
            or145 = or143 ^ or144;
            or146 = or139[0:0];
            or147 = or139[1:1];
            or148 = {or147, or146};
            or149 = or148[0:0];
            or150 = or148[1:1];
            or151 = or149 & or150;
            or152 = ol17;
            or152[0:0] = or145;
            or153 = or152;
            or153[1:1] = or151;
            or154 = or153[0:0];
            or155 = or153[1:1];
            or156 = {or155, or136};
            or157 = or156[1:1];
            or158 = or156[0:0];
            or159 = or157 | or158;
            or160 = ol18;
            or160[0:0] = or154;
            or161 = or160;
            or161[1:1] = or159;
            or162 = or161[0:0];
            or163 = or161[1:1];
            or164 = or1[3:0];
            or165 = or164[1:1];
            or166 = or1[7:4];
            or167 = or166[1:1];
            or168 = ol19;
            or168[0:0] = or165;
            or169 = or168;
            or169[1:1] = or167;
            or170 = or169;
            or170[2:2] = or163;
            or171 = or170[0:0];
            or172 = or170[1:1];
            or173 = ol20;
            or173[0:0] = or171;
            or174 = or173;
            or174[1:1] = or172;
            or175 = or174[0:0];
            or176 = or174[1:1];
            or177 = {or176, or175};
            or178 = or177[0:0];
            or179 = or177[1:1];
            or180 = or178 ^ or179;
            or181 = or174[0:0];
            or182 = or174[1:1];
            or183 = {or182, or181};
            or184 = or183[0:0];
            or185 = or183[1:1];
            or186 = or184 & or185;
            or187 = ol21;
            or187[0:0] = or180;
            or188 = or187;
            or188[1:1] = or186;
            or189 = or188[0:0];
            or190 = or188[1:1];
            or191 = or170[2:2];
            or192 = ol22;
            or192[0:0] = or191;
            or193 = or192;
            or193[1:1] = or189;
            or194 = or193[0:0];
            or195 = or193[1:1];
            or196 = {or195, or194};
            or197 = or196[0:0];
            or198 = or196[1:1];
            or199 = or197 ^ or198;
            or200 = or193[0:0];
            or201 = or193[1:1];
            or202 = {or201, or200};
            or203 = or202[0:0];
            or204 = or202[1:1];
            or205 = or203 & or204;
            or206 = ol23;
            or206[0:0] = or199;
            or207 = or206;
            or207[1:1] = or205;
            or208 = or207[0:0];
            or209 = or207[1:1];
            or210 = {or209, or190};
            or211 = or210[1:1];
            or212 = or210[0:0];
            or213 = or211 | or212;
            or214 = ol24;
            or214[0:0] = or208;
            or215 = or214;
            or215[1:1] = or213;
            or216 = or215[0:0];
            or217 = or215[1:1];
            or218 = {or54, or108, or162, or216, or217};
            kernel_adder_4bit = or218;
         end
   endfunction
endmodule
