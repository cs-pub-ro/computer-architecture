module mux(
// TODO: add inputs o_w_out,i_w_in,i_w_sel
);
// TODO: implement mux x:1
endmodule