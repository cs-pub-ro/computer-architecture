module fsm(
    output wire o_w_out,   // found output: 0 - not found, 1 - found
    input wire [1:0] i_w_in,    // char input: 0 - 'a', 1 - 'b', 2 - 'c'
    input wire i_w_clk,   // clock input
    input wire i_w_reset  // reset input
);
    
    
endmodule

