module alu(
    output wire [3:0] o_w_out,
    input wire [3:0] i_w_op1,
    input wire [3:0] i_w_op2,
    input wire [1:0 ] i_w_sel
);
    
    //TODO: Implement the digital logic for the 7-segment display

endmodule